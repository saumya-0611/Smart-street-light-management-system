PK   ���X����.  `_    cirkitFile.json�}�n$7��44X`Pjx�$���3�c��6�93�6
yu��J[*���h_�<�!3KRU�̊���z1ݘq��d����^��]l˟ڛU�ٶ�����zss��ˋ���<�-���]߬v�Տ�������������6��m�TWgU	[�V������&+�gL���Z��Wl�.^����|	-��8V[	4���hX	l����J�1`%�U�ƀ��VV[4���N�S�z��vs���V�.��(X��2%
�����Ȃ�\��<��^.���de��Rd�.�̖]���ҭ��.X�|���x��Ph���x��P��4Z�C�7ӽ� �%7���"�Z@~~�@�p(�CZ�C�,�"
�G���I��F�p(�-¡ p��[�-7Z�C���h�Nx5]aE˫:+D�3�:��JWYe���M�qӢ]���YW�R�2S�v>��Oe�*+�,j�����S	��F�p(��S����D]g�-�2ŵ�Ĵ��U]�ZkY�Bf���=Z�C�7�������6ۖ�k�$��vs]n׻_]�D��
Q��Vg�`��VT�MQ�U�Uە�cw����D��p�NZ�YU6YW	�TY�,:�UmÚ��X1��($�Np*����m$��Cl��F�,�r�8R����ư��y�)�lV2��1��xc�C2��|���Z+��8�Z�5����#qi����c9��0~NO�V�֊���!���+tm8�3٩2S�s�*���-�<o���M�6}�V�V�����3̜���*�U{N�vRt�[��+huG��Ӣc+C�;C�;Rt�[YZ�YZݑ������8i8ȉ�qb|~�X�Q&)>N��/;�/�_��K^����ߍ�JS�~N��u�f%戴1^J-��yV~1�+∊�F�'�痉��G������
5����Z|��_'�q�B�������(����.��l�Δ�۬*��8˝u�Ei�=�ȉ�����䑨�8��AHqvSbg�h?�G>�*�p��K��x_�U�L�:�+2�k�U�4����U'�J�uϘ'�q��;[U�i=�O�[u�UO�������&#b��i��81>�=�Xı->N��o�"�q�E����[҈�Gk�������6b��Z��81>�!�X�->N���$��
->N���d$�q�⋹ޠ���}ӟ6s��x�������3����Ϭ>ޏ>{�)n��(C �tH���f"o�Y}��{fu��W���]�s��!;Rp�on}dW���U`Z���S�^�"Mptmn}dw��:��Q���0��XmЩf��HWt�r��j�ZP��ƽ�ÃcWs돏�έ�cJu��F��ǸW�z8h�����жQԫe�8��](ԻS��n�x7���K�� ^͑�xE`���bL�X̫q�G ��G�=�h�0�a0��6�x���U�8�؆i��j����� ]#;��n��t�@��1$�z��UO����� T=흂��AP�t�>>H>�z:�������X}$o'�>��&�
ʔ��71�NE��w#I?1��_��'���ł�CA������ه&f`���bvV�� ����Hd�;v#�'���X��?��D�O"�'���i����L1($�� KI27�V5Csr���yur��
��P�ޞ���.�_L��p��p�b��SS#���OM�W�0���a�mqLO}7p-�ݩW������{`7��IMA�ޞ�Y��M��6�M���tm]e����u����E�[�L̕���}��S4-�t���}c2[k�>�t�zu��f����箅e��De��T:3�2Ә���sUM�T=��κ�E�ʼ��r��۬.U]Y�I�_P@TO���FH��i�u��w����Q�)Ti5�vP���������z��߿p�������d"A�m4���w3� "���@��HPo""A�-4���w:� "���@��HP�""A���$c��!��c�AZH2�M%i������d��J�p&2��Ɍ� �r�7WHLd�{�D��̀SIn^ �Df�9���4��@��H�pG�cIf����4��@��̎2;N%i�ہ�.z�[i&s���{I��9���4��@��̎2;N%i�p�SB�������J�^���ŗ
#5��kx��^�?h�:��A�5���F�!V<�Kh�:�B��+Ek-�5̿O��yBh���0�>�ƙCȥځ%��Y�i�:�(B��q^�X)��X���R	���0o>��Hȥ�u	�aN}�3��K%��X�|�4g,!�J��%������0��K,�6���H	a C-�R�K����'R��L$�?��	�"h)|� >�n��h"����R�v� ,ȖO��eB�E�FR�Ӌ���h#y����L d�'R�2��"h#WM�.�E�R����2Y�'�f&q����DJX&(r�)a��,��d]a��,�tO���R�"h#����R�v��l�����b)u�В�h#i���R�v��l�����b)u�L\���u �b)u�L\���U�b)u�L\���5�b)u�L\����b)u�L\�����b)u�%� hg�SN�����DJb��ܤY$RT��fJ���y���.�R�~g�k�R8cy����[;�uD�ao��\14��Zu]����ٟ�ҝ�14N�A��N�w˖��È�a�p8�f8O�#h�а8u����b�,�:�1�'0��ch�X1r�ŭ�K�ӳ�:��6.��}���9קGoh��iO��|���I˧��p|����§���{���)����m{�_CgO4���AVO�Mh�j)'Ghk)'OhNk)']+h�k)�s|��]H9��_S�����pJ�����zz�'���(	�8Ma;iX�:mFj
14,>�sSS��aq�|�	�)�аXҰXҰX9$4,�4,�4,�4,�4,�'Y�~}"f�><�NO��AHOO�AsA�Rf���<=cM�K2?��4h��XN������@�����OG<��Yx�A�O�ihr_)��r4_�4h������@�I,�\�RNb�f�%�r4�/��C,OY�v�%��{�����!������ "4d�%AD$h��K��HА����!�/	""AC�_DD����$��YI	��� "���Kc"�6��&�ۜ�pSI�g���Df�9�񦒴��K���~s2N%i�����dF�J�>�/&2;.��8��}�_Lt�7�Nf�������K��̎2;N%i����dv�J�>�/&2;.��xJA�_j��	 �����RɰF��RK%��X#YI4��J��%�F���h 82L-�P�K`�d�%�@p\�Z*�^����K���0�TB�.�5���D�1aj��z]k$�/��#��R	���H�_ǃ���u	����$�SK%��X#Yi<�e�0�.��Lȵ�X�_r���](�Z&�
�蒋���2��"hcY��R�v��k�����b)u�L��X�_r���]&[m,�/�XJ�.�-�6���\,�n�	�A��K.�R�˄d���e�%K��e²E�Ʋ����\YX&.[m,�/�XJ�.�-�6���\,�nZ[&.�蒋���2q�"hcY��R�v��l�����b)u�L\��X�_r���]&.[m,�/�XJ�.�-�6���\,�n���A��K.�R���e �gd��KI��>#�/^Jb��Y�R{���������{F�_�����s����ao��9Y	��8u:Ꜭ�bh8�:6tN�_�G���y�s����aq��9Y	�а8u㜬�bhX,iX,O���/�������r��Y'����⥜�"p��I)ିx)'���wR
8�/^
��#
8�/^�ɖg��K99(���⥜��Y	�K�H��x�_14��tt ��K ��§�x�_14,>�����a��� ���@�OG�bhX|::�g�%C�bI�аXҰXҰXҰXҰX�d18�/^���	��/�$��Y�RN���/�t�����r�XA��⥜�����B��d?g�������rھ@��⥜�G90�/^�i�����r8�/^�!��/�?٭���f�Z7�\��������[�^�u۬�7�Ͷi��߽C����G�j�<�&C���1H�؁(�f�A&ݧ���������'��΃�S����b�F���%($�A2>U�iT�
�a��D2>����~D�4�ލ�"5�n�*�j� ���hPy�(�N�+�8�3��eM�-N{��2a^-q��0�F�g0o8yE�My�ɕ$ge�O�8̈́z�ȓ�l2�vE@j����^>�gI�!д����*�Y�9I�g��I���<�~�q6�<�V����ޥ�1>�4ݨ�� ���.�v�b؈z�I���L��)͸�Q�ɰ��Y�w����u����sT����<�n������Z��̡��1����p��j�k�y��W?��^�m?n~j�Uy���.�9��0�ߟ�B�zrYd�����Q/�D}Zk%$ �\2�lӗX9��(=�O�	��";x���UD��3��yV{ `}&!���O�s����%֤^���KS��^d�
��z�j�ўc�
� �l�G@�z�D���h�\ka� �kIlzh}���i���Π�ˬ8�~�ә�ZD#�zGJ<�D�#�3�X4�Wɴ�\�uE���bΘ�tw�ivyE�V���IE=�jq:Zz���Z^d�#�H�BG���/ˣ��>E��_v 95��L��ly�5�jy�����e6Q�環{)����b���H����s�+|�-��_����v��c����v�ۍ�������~}�Y���]{����M��W���~�\�����s�+�Ȅ��s�Hh�?_�D�����Hh�O�D���tqHh�O7�D���tuHh�Ow�D���ty��@���i�L+^��aqXWN`^�2ؐO����r���5�Ά�XX����`C�E,;�	1^r>bq�e�!i$�y#������e�!m%���/��3�8<Z1�	+"�P͆ĞXmX[A`m{��a��H_�6�*��d�Ov�F�
�i�ӑ'лщJ�����"ّ6��b�eQp���p�n�!DR/�Yv�� ev�SN�ٖ��>�{Jp��.�c���!\������#����]�G_.�E�3�I�����K2�$��G�NZ|�[����#�-����{��`���'��V�}�t�H�G������
䴁�Fȩ��j�G?�95Bv�c�F�A���d�0&D8
�q�d8mh��rj�~u�Z���1BN��/�Q�:f!Fȩ�uGjR*�95�0yD0��t|,�F���1��d4�����d41��H^���|���c��ёk	�S@h�
�'D8� v�:��!��y�rj���T!��Cb��AJ�'S�8�:�!Fȩ�=)�:��q�rj�~?��cb�����C�C��!�F�w*Q�:�!Fȩ��s�4:�^�!F��2u3>��� �h6 �P}���x��������-�sS0"��m�U�aNK[Lg������|&�^�s.��l��5<�3W ���#1���)�i�a�O��?b<�"���ߘ�: �Iٟ���t���H�9���A���C^�S*A&`Va-F^�q��"r>cUdHy���)�f��6/0���z��d��KH�3�@���xz������[9g'��v`��E��iǦg�g焁Z`���=䳯Q�>O07wSڦ��O�n�����Ġ�?����O��������_�(�Y��� S�L ��S�����:���aI:}@3�M﷛+K����\hË��T@���SL ���Q���3<I;w �2Qb�(�> ���D�e��2Qb�('���b���;(������S�����0{�t2����SQ�����#fg*���O�嚝�:-�oc:���\��IA�͍�a��O'��)nb\ ^n	](�9oJ%D�k[;f�"+u]e"/eQ�VUU$�����dˍ)��e�i��1����Ta:ו:[K3�~P����y�e��Ce���T:3�2Ә�ю�\US�՟xg���Z��ު)�)���RՕ՝d�3L����)]�9��N�A/�Wt�S����z?�����//���P�	��U!����]�q��zOf�]}�Å�h���G"?��ӝ}�և��^?+�ϖ�s\� �]�`�����-|o��$j�pԇL�,e?{��j�3��ֿ��,�1|W	2T���� �cA%���+���}M���C�5�V��א��4} ܝ�t����SEW�U���G C�Q�0�x��?z�B<���`�*@��Q�Md��������}�q�
�x��������^���ڬm���t�Vv&˻�X^V��CI�W���:+�\��ϝ�S]k�K+�d��c�7��t�*3������hÚ�����v�ۖ�vZJ�s��5in����^fQk��.kl�eʸ�;v�0(nx� 7���7u����w�����*]�,�����~p��~��7����P�x=!�Ǡ6W�oI	�q8���pyUz F&��ȵ�:}����v|ay 6G�]��� l�h����< g�^��� �Ũ����18�2�/r�w�.e���Z� N�?����-~�ˬp
��b� \ʚ=�����z�˜4)s�;�����z�K�p���L�x������J��g��4�����u�g�����O2@�1�or3��.T|��(�\WJ��e�-�%���0@����:� *��^�7F#Q�9�+�4�@�9��ФƔg��/@�rK�嚿 M�">˕Os�����꺬�k?e9��~��v��w�����Gb�H�������#>�����Q�T�����	��#<����o��~4�h~5�j~v�����g�ï�_���������'��8E�S<�!N��E<�!���v�a��:��ᙈp�g���D�:�j�Z<�Z�����僪e�j��2�L>�L�*��(l"��������y��7�fu���y�S�"/�Jg��O5&�E�ܔ�tM�J�l�'���/���37������Wm];�g���W�a[�7���h�����\�B�A��S��޷�ܨ+e���UVأ��vu�v�~m8���������������_}��ܶ�ݺ�W�?������vMt�ۮo�4�M����^^�T^�����M�{��߬�������޼qr/^w^���]����n]]���۶�y�޶����G����}Wֻ�m��pX� �p,�Q��z���Np{U��*r�N���J_��0�g��h�k�Z��+'�BȦҊɬЎ��rC[�D��J���P���Ǧ�{���_�//�7w����첸��l�NJ9���i[���u�o�wNΕ-��@��8��B�p�T��I�<����%�T̂�I�&%����4�I30i�X�N�S���q��uT*W��9�X�fA�I&M¤i��<7W���RZ�J�� �R!wc�B��J�̍�
�+�m�X��A�~L��E.����i�����Ǌ���_������_\��X7�ol��M�eƸ�!T�B��	̊�n��4��m_����z�����x��P�)����\��o��{]\�Ś��.
�L������x��������T�k �п�˅T�l�c��nn�w�u�"c�u�;�ee)�����uj�l����n�k���:��ߞ��͇�us �4��]���UR��A��W��k�pk;Rśr����޶7Rr�TU�4�?�\�or�3am�ۜY��)o�7w�!YJ3l��S�a.�t�NH�`2�0��;���myӴ������������gu3|�����O���7���a�oXr����v�E�lۻ����/����[_�r]���V�Nu�VuQ:���V�&��s���Z�$Xm�cJ�e�i
�"�y�U�fZ�F�Lˢ3�v÷cF�Z�喎[�)�κ�*��˓�U�u^T�s�]�V:���U��)+k��&X=����ͺyu���o��?^����ͫW��+��W�n�ÓW����|�ۼ��߼�8��+�����W/�z����X�o"b��m[�����Ca��������Q�~�./��O�v��s��ѐ���.
�R�z?������f�yt�.�����4��ص,��b��B^:f\�N��{��У�L���γ�i\���uSoz�Vi�UV}�yڣm|{������4N����+{�G9�]X�x��:xMj�B
Ί�2�n�J����%h?0�;��k2���>���Ɯ�O=1E��2�����D�^-�pv���"�������W���qnȞi�5+\�ۢf�ȧx�U�k��.���d�W��P��Ǎ�|���c��� c�e\�L2.�~P��85|��_�z�)uЕ��\��TA�-�4��̚���������fV�������|����_�g+�R���kQ!��?�C&z�����W%��k�8�5�mڼm���Q)��� 3h�ME��e"��3o�x���dƁ6�3�rހ�X�l���:�x)��?���.���q�U��t�D�<"G�>�c	r$G���:<rr�rz�0E7�+�soo���ڗy~��LSȧ�8ٵ�u#X���8;��ת`�s��0�v��=Hk�d�>ř��FԶd����Q>����Q`H�h�DC�ȢЙO =�pٹ��X-�>Ǝ?��3�2Ea�3�����t��5N�z��>��t���/�c�֙��e��֔9����T1��� �Jׯ�F�r���F�ɛ,� т�N�,(�%�Z
�D��U8�-�Gf��T�JT�~�,(�T��J,�-�e�HJ�%x5<����I�OF���b<�D�:<�txc��D'��:&UG�T5�w{z"�uƎ�ӓ<Y�H։�}�$��}`t�'ڌg9�ߵw��R�����{��.�A�'�T���������C�/�|Ͼ������g����[+��4nT�~���6��v��A�;3{DO�� ��cȭ>���W�����_�O������#�7��&�K��7��v��m���򦹛�7.{����tN��#���|Ìc�PV\���:ȣ��u��γ�,e�T[dZ�1��S��M�{5��#PB��H�]��!����?���΂<�}���V�������J|q�skB*���U�b�2k�&��U��'�{2��g��ܸ0��fަL���R�+%.L��̊eL;(��Ɯ�ٜ?�����g��K�ز�в/�{PB�3y3�R/m��g��-�W��V8�BH.���/�{P^.�-/�i���OF}@��o�Џ����C��z����_|���߾���7o����o����o��h%���qك7=���]�ٿ��ߚ\�w��z}�桝�]��X�>|����>�������vsӼ�\oW�����<)�]�g������-��/�����k��x�/�����*Ө�������Q���
vRZR��7�{�#���i��7�{7���E��q^���e�su���N΅�;:��\��U��kim����Z#��we�lC.�e����M������د�{���??���쟺p�\0Ʉr��
�WV1���o�>��z'(��'�;�����w>g�,���Z��0ô�s�;�+!|>TUxwx��	J�iu�/?��;�����\1�׺p2/.���ΝO[����t��&(M�'�7?�����M�\W�ZK�H����$�ܸ�3w!�2����_���]�s�|ή�C�+��Ѕp��RW�Q*�:�9�[���	����o�����z�_�?�{�k���3��O�0Y���F��o�,\eFr��"�6_�{�n �wO����V�6��.�ͯ��o�~����;�^����~^7�^�v��{�ޡ������o%΢9����2���������6_>���v��v��}����.���o>7�cZ����ϱ>!�������}
��o89�4Q�Oz�����)�:y^��f��Z���������>����[����R��߾~��{��ɬ��Y_�2RJ:�G	�?,�������??��\�/%�v��?����w��crc��RQ�P/E�Gb�I��v.	�Ix\*E�B@H8*����K�`k~���"I���Te����������4ے��f��g��Iţ�]I*�J�d`�&��1}@�8���.�8�X���i��Rq.��a�Z����+89g`%��q�3�:nH5=V�\=�ػ�H)=�脌�H�I-�i��2V�̫�^�Fk.fyY$�)�����Gr)�Zf����Hlq�@1*��A�kjwƄ FS�v� ic���������;����'�{Tj��vS#is�3��P	[;�vn�>:D���ǥd�	ԣ�P)h(;�8�[4i�9�93�Rډܹv��'��q�)��HV
J�2fZ�Y9ŝ'Y��R��A�	���o&9�����̓��d\]�<��K�O�ؑ� �:N��4����i��KNJ��ً�M��)tb��<|s'Ӭ>I�Q�9� 
�K��HS((F��®&h��~���l�\�ǌ�
��+f�ٌ���V�7576��E�ss��=.���p1�'�b03�u�f�r��Sk�M���x��'�ς7w��ڜ�83*�A�SMBK	�b��y���x2x�rV��e��K�RLwҒ2|j}&��W%�����e��O)��Iq��_�:��|�3J	-�Z�)���fwP��̓49�2�[�f@%��[����$�����ey��*��~?��"�*���*?�Q�C]f��LG5�;�w��Ƅ��`9�3��Y�t��g����e�Xi&y}p+�y-l�r�9;E�'t��}��߃Q���ς:��9d�H����
�����ŀ�7�;�"��ddv���3�瓊�S�����	��x�Z_38�DA�xsW.�15is3���ܝ���p(�B�S�cT���qold`����	
h&s��2X�
�\gI'��3I`���AsKAI0+��\A<i/��f`��v����f�h�B�hȞ��JE��6��;(�r

�F���͉=D�x��oɐÍ��cV�x'��_(id`K�A1`̱N̨�(С� �
8�f`��(�d�r�⸐�O�d�F-؆��c^g��6˟�r��o����ŻܞSj>����S��I��ht6�:��F7�7��ʤ�"�W�@���hc>�T8�=�`gLA.-9���Lg��mZ ��rо���*�T9 ,5�e���s[������� �����e��2�e��;�T<4S��jTLķr����J���	#� l�0�a9��3�;nj(q aT��h��cC+�
 ��Y��E�L��$�D�IKje��;g�C��6��F�LzV�)��{Ge.�[WA��ȧpC�S�KyU���&�ŀ�$�8�{���Qlgg`#3��M�������d*J��[j���֐-��R/fa�9h���2�G���ZF	��d%�2�J=OV��������Q�P))�ֳ����R�EPz�O�/�\Z�&���ĳ��%?�����@���QZ��"����h��D�����;E�q��}V�������ݮ�뻋׾?��?���m�Z�ܗ�_n>~�k?��&�����������O�]�]��r^���PK   �{�X@��)  /   images/0931d3d0-b3b5-4a2f-bea7-013f7f069bf2.png�{eWM�5��I�� ��w�;�a��]�kpww'@���;�>0�溟?�~��յ�ԪSGj���Qj_�q�(�p�|�@@@"  �`��롭���w�t��熀����1��
W�,��sރ�ch�!��թb���A&��A怳�>���P1��c4�{?�ԗ̈́�p�i�7�o���q��'Tj��7��+ ��x�t��5��@�4ic����}���R�&�%��_�&D�]���]f3�d�Z��4�����H�Dc��K�j���]tЋ���2������o'*�k7}���������vF��*���g�u�ҴR��FR�(��y�J.���{���>u-y)��ȕ̚���7���/��L�B^��Yz�v���~rm�$�=ھx���%����$�p�(�ێ)�b�d����RW��#|t�#ge������&$5O�v}͎��l�<��էa```v:_��(�m�Xd��!�wgKG�}p�9��q��Z����*��Qp�!S��r0���t{�M�����/*��s�OV���1����3�eȃ0 C1�H�1��Z/[,V��c���~h�~��y�o���}��!V0oڦ���\�#�<��n�����E�v4̥]���<@ �!T���x�ف&dlJà�m������b���-�Ɨ��u�(#x��)���Ŗ��7|x�Z�j�S��(u�2hU����Y��W������ݦ���Ԁ@��Ga߾�X�Qm^�{0xy���pg����w�ל���/[��cu<َi+�u"��ʨ���۳��I�#�Uc�&�[������׉������ܱr����X�rAĈw!��/��6I�˻/Ty�O�R�0�,�8*ɽM*�}�վ���?�kV4ʷ�%�Û��1��[��/uzM�g�P��_a�'y�|�1���!�cQ/ے��恑�x���w��0y���#j^�gX��n�DT}ҨL�@�"9�=H�y_`�~/*�W%�L�kH�3DB�5,�W�@?{���<��������ѻ��껀��	��/b[;��W.�܍d~UI�o�/����R��6�P�wWа,����T�^Nw�A�֪�����%����t��'7��Iy�-�r�|��cC>�܁�������k�8TZh%嘙�k�,lV3�U��{��T��}@���旜�4ӏo��g�.��Bv���sfK=s��:����ʷ���L�1����]�j���1� ��6��uj�[~|�eĔE ���^���/�O~�бd��v�z�7s�2��L��xm�$dr~�t��������L��E4O���q�~�k�9�C$�@«��
0*�9�A-p����"���A�ݻ�ޜ��۟�6�[t�s~U��q��x���}Xń��y��m2ß���É���R����[�gb$Q3�AȆb���$l��TDl��4�m���NIͰ$��te��S	�)��>�9�'���B�Ѐ��k���vgCFt-*�P�ط?eg�Y�ny���N~�
�57{zz=���a�	�ãNݧq:.�"G���-D���e��'7u�\aww���jk㷎wuj,8˚3�"�/?*K��:�%�����v�v2�1�bf(1?���4.�I"ɍǬ��^��k�N���ɢ������"�ථ�T01�Ѝ=�ꊟ��:&2��f~��P�O�Lq�?���N���r��`l�e��ܫI8�������)�,����_��K����>J��r�9Ih~yC���)!���5�н}������[����T�'�-�>*0��ʏwLx�� ���8?�|��PK��O)�I/W.�v�x;�0p�R�l˘�)ո|��,���/��'��:,�d��T������u�b��
��%Br���w?���iI��Q_bu���qՑ\�#���#��(a�t��qeg�� z��"H����l�D���b���.�ө�n��\{[A����a	{Iq&��K�vGm��c��q�h9���
j�h]��<)Iw��q�U����դ�倛j��^ ���������\���D���->�ao��'e�讛���K#��L�FPJ�p���/�_"K0v��5���h�	�80�kw��t�y�V�����U���O�Gl��t4�ʱp�ll?%�!7,5:���n�(�6�,:��F�~��%��OVfJ�z����I��P!�����'�A��F�3���촗��p�(�?T�E݅аA�F��snA�
�ϥ�=�̴�#�b�gV�-�g8����;��'*.U{q��  4E�~���N�I'���P�x��A`�*p���C���Kښ�'��O��A�/6���ކ�5�-'_dD�ۦF����Ά�()��]�KLjQ�E�~NMq* @��5���C][���pQO^x�/�-�&y	��� ���e�lYfʷ�iߝ~�k����}�6z�{t����͞ �N�qC��:;1���ަ0��)�U���vi��C�s���W�C��e�C�t�4��zp�X�_��W�����|�C���Y�å��h,q�W>x����q�������Q���Q%|u� �� �!lg]���i:���x��0�2�p��Trchuy����^@�xiy�+�Aa�N��7���]@4F�&�e��Wl��ȶvu��4��J<�_�a�n���^����h�3� V�ɏ�0����f�N���;��iu�K;~���j�۱�
���	�p�9�����Ew�'11���>{�� ����Xi��n�^^���H��3�@� `���п�jYY(��A�tޠ�������S/�:c��a�l�z9�51��ǡ	���.�ɘ23��K��~�h����~<۹��c`��.-0�`�2B��Ť��M MH�c��2�동k=��y��4ع޻Q�S &&�0����f�~�Dp79y���b�2��L<~�/״���Wz\y�-VSYؓ p��y�5�m��(�uq���{��1��c�ɓ��Oԝ��CK� �4�q�j���Jt�ru��e��c�^�Ӗ��󅤋)�����iP�rp��������Ѱ��K��9��L�����l�J��,����@j�z؀�8��)�����:����P�@��Y��+�;���?��1�p�F_�ϟX����s������>s!;�K�.��?&F2[�i&%�,ߧ��AE�o��U���n'8���?.pr|��~��"�9������Be��t�0��Is��^-�����V�k��]�������~�2����ԗ�\���I�p��Ʋ���0�_g���)�t����N��SR��O�A�O���� �A�酵B)o�&	\��ᖨ�q���?CK)f �����}�Tz�������-wfm�J�ʯ��&T{Y3�E�\r����8[�O�����:L\�A��.�
2���N�;&�i�Ut�����s�e���K��C�
B	W����n���~��NM%�����Δ	[��]DG(9��(Hs0|��T��a>����{L�d���H�ю+�S���ʅ�'$X���P��k�ζ�iS6�huI9g�TݓKև�=�w��$�o����''� �;̽��������q������أ��}�GnȨ�D���Eϭ�z$�mv��C�C�e��a.���}�î�d�"��_:|�y�,4gZ�L�1ɺ�z7P,�eT�_��h�Y��;u=�A4u�U��A����8agF��!�@�� ~7[��k!߷Qg����÷�Da?)�%�UZ���=2X��=o�5�r�+�j3y����s�$Ʈ�}��������*9��2�p�[i����~m�(���n�g��Y��v����h�T�ɔibu�3�T=}�"�MZ�:-6m�_�>G����Ↄ1�C�����Wwt�I���i��f	F��P��8��7��!z�Q��Y䖫*K�_)��z�C�r�;j��v�-�%�%�XNi=�a�[����x��Dww�Ϛ�h����Jj���hQZ�;�|����ܭY��f�
=y�ne����ֽ���X&t������.���t�@ � ,�˂�s�}M8Y���!�� �2"��>���
]��b��@�16����iE���fO��Zz��61�Dg\F��,�N@� ��)舞J�����Mm�O}ɟ�C�`�}�!�7���5it �dC�lL�$�I�@0*`Z9��2��`�x���bM�=9��m��:��?���N�X��u����Q����;�#�ï[�~#Hqi�(�O��P�w���w�����"	���W8�@P�&�u�kg���J���;�z3����{'�&.�����zT^����l2�>M����!UG7>�o_�{��r�&w��/6Ey��~��<kB���׻�N�I�p���f
�&u������C�Ǧ�;����U�1�������iDJ$�w���v!sT;K�=Տ{r���Gj�{hN����q$���ͯ��X#)aG��Gy�^��	�4 �C�	�^�X�&1�O�֫����D)�Fg����S�L!G}���ϼ(nq9�2�tR�+��eF���#؉ey>�NR��g��?��tBy�L�}�Or�:\K��t&�,GY?M[q+1�R'S�Μ�4�G�oֶ`���3����|���d�H!E�BΛ	��.������W�ɪ���!}{q?ڃ{�fl�|�J΁���e�8�ސ��ìs}J_n��R��.���ι�7r/쮎}o���=���0��B4	�
κ��ez�Pބ�O+��MMf�һ����I��3��O6����L�?fn&�ٹ�I&�)�z����= �w;zm�)�'��'|�����\���~ݚ��������>�� �=����L�o��ę�r��{�#½�o�wm�?^���]�s-7��0�B�����$���\�D�O�c������&yG˓���43�6Fcq��dUK�:4����Z�X���(��A����wā���#H2��BLΔ� �u~� .N9w������o�^�u2i�x�5�5��w��<ay4�˳HI�/��y��X�׏�II�D,���Hė�>����S�����S�_䬺i_��'a�e׎3��f�֫G	�?Kо0l$�2�4��,���wItN��f��s]w�=ےqh����o��x�@�|Q2CX0��*o(��r_^Q��ֶ����2vf�=�6hu�B�M���U��;=���s���~	��z8�B��sJ��W��w�Db%�������{��2m�ݗK��w���R����&Q,����U�UL^|�Z�$�%���d�GҫwIC���.����~u=2jc-�e-�U"�mo���9����}?�Y5��8�K��~��b��(dk���#&؉�A2+��4�2��&�(p#�u���^b��}Vt=9�M�q;�u�����S4�9X���N�A�ӗ��(x,'�.��r�j���n�\��K�MI�T�W��2�����u��uP�l�����ّl	K���a҄X� Oc%%�Ж3���J�Sd����R��Yp0�0�tXF����0E�Z�T����� ���#-�B-F�܆�?�]�<�K����o�	�$-3</M�_�N�f̊��~�x��)�Q�En��k���?ĥ9�ZY����x����Ìi�{��d�W2O&E��_���'*�N�
6�+<�.R���S�^�G͊o&BT�7���3K�����ݍ�o�0~�0���Vd���48B�Df8����ƾ��Ѻ�ʑ|r~'�"Bm����wK�lN��b�-�37��:�������h:`h�t�2}���;��-�)
6}h5���LY�� ̓^Mj{����6}�:韬�sX��е���'�W�P�g
�l��LI��g"�P<A�9�a#�w�S|��1�H�8@_�����fP��qQB<��6��
��T��I�as��!S�����S#l��}�t������P�a�蔏���un�(-@��{XV�J�@="��u9�f��6]�8c�π�n�1mڒ����d]�^�h��c�M�֤�8�f y��} ��Q	���x�^�;۸���L��ܢ��:f�$/�駭��B��,��/!��g�cۓ7���:	�%~ �J�O?��������X�sG�</W��Š���f"�
�u�t�fC�s�������4�;tڇ	�c���;B�dF��3F��
s�U���o�KE}�|�	=��9�&�Hs��|�C)���	c��*�n^� �S�y6A��/$=�N�1&K��i0�h����ߩQ��L�\�%ޑ�I�u+'���U�U���/�A/3� :Z�AY#C�{��:M%�5�-�2���h`���B���fϩ,�f�K�� Dc���	W�@'B$7i���#�yDh��IoFb�&��_B�����4�� �#�\c�aA.�%��ھn޷��UjU	,C��^��=��EU�($bP��rq�℈�?���BT�Mm�)�Gj�d��z�㦨�OzG��|��U�}�т� �.����������wb���ٙC,ddD$�hQ���q#�� :�9�1=#�Ȑ�X��Ǵűo����B����v�X����S%S��!�g�VrLo9��/��:}s���~�<���j��h�`D=W�g�������|~\��<va���|?�=�ď��٬<
?�vJ���M�C�
%�� �T�h���>�7~�*�į����ȵ�H($�
�Zn���E��v��g[�?Ĥ:¥L{�Af�b%*�����3T������G�i
ߘ�jih���&��xY�O��fB�,	n*�×}��?��V��NeV̛ X�)�S�';*:�2<8B���:&5��їf+�N����=�V���2��/�)~Չo�u�&��N���v�y*�'����&����޽�\}��O��3�ןf]@��o�VA@�<P��]�:P��1W=���k
9�����5�o���~���b��J������qpW^�W����q3D��GX�a
���9����������d�o�S-|�>KU�@/�J�t���������x��
����shu��}�h���_�����|fv��o�M���I�>SD�K��/]�P|w��=�	7U�2��mv���٢�I�D~���z}��	����g̻�a�&zF�#u�F:��Ʀ�<CHJ�����m�{�|Э��Y�f10z��W+��C�]�Qz@R'a��]/	Q�O�����Gv�k�L~�x�Jn��ʻ�[��y���bI��H�lۗ�8)ώFnE�P�U�[cW��q�y�t��S��9�"�
|X��:[��J�������O�4���d�m�7�q\K�,"y�=�T��	C��'��c�J��ʕ$�&���į��#����1#X����p�E�.Mw].�K����1���	@���87�N�'Lw!6�ۀ�5���=�?D	��F�~�	ن�y���<9f[T�	1+�b+8�m�R�JO��Ũµ��Bgw��?�F*�.\��$�x_#���7��;Yn3�j'�����=]&϶��D��ID�x��>k�7�_c |af*PF!@7S�� @��o��]}i��f?�"x4�IwA7�{y���nwȆ�4�> �.Io�&�p���kަӢ�֌2VبXݘM����X qJ������Z��=1���q/g*0{YY����;��d<�/�����_R���*�[��Vݤ�*�ڜ�fS��O�ʲ1�)N�CɎ�'�������5�bc�s��ID�Ή	�N�u�\����7S�kM�"&\��2ԥ�^:�s��b�#�po"�V'-#������Xkz��^>������FR��Ν&��v� Ix7���^�Cf�� �H����|{�	�Ce2&�?��׵��l9�^"~��o7���C���/K��~O�w�&G/��qvm��(�&uv����7{��Y|3n<�#�Ɂ�Kl������v�X���(��{��!0�2qƪ��\�C��D	f�n��_4����Gx���^&���|"�V�-�N�����/1v}ŕ�����oӉk�]Z�4����_��t�}J&��MP�G�h�	�+��4O����Zy��m����[�^�RXi7kz9��\$v��V-�>�_������Λhp(��:;�{9q]sl��wy���x�	q}���EGA��+Sͫ͒D����A�Y��oG��G5T��E�]-��D�ep/CX�H�QY6��0�ة��hK$���J��N�Ã�C��k7���ON@���,2����l�r�����p-�'J�\���9�����a��e.
B5I���â�s����.*����=�K�?��4�f;�:�׀��B��B�aJ����1V�O�)��/�E��Fmcڟ��}��_��t�l�2��.����1��g������6R�������lN2,8�
�]�S�����S�}U�@X��Ɔ�Mve;��a�0
$��P)}��7#.�T��G\��lp]	>����%t.����V���΍%+[J� �D��h�li��z�X�� nw?�x@%�>JY�x��h�VP��l�Sw~Eji��u����|�M�6���j�^�n�JH�ؿ��dbMߋ�̬�����F��U�!�k\��O	˴�͌7T����r&�m10ͬ�:�j�����ז3fU��Ѳ��W����������E HRBt�U�(�}f!�JBN�,km΂L���HVӦxG 8t���h:�A� /ɒODO;���;�zo�;".�G�,W����%�D:�C1C�5Ŀ@������z)�Ɍ�#�2���OR*dҞ:����ıd�b����t�q���c�׏��q�s�{��RQ��+�ж�mi��s	�l!���UͿ�!�
���)�;�;��Y
c�)�PCp��N�G�_�E;Wh�̲e��	���̲f���56�eV%���e1�~숆�գ��[�+�������R��h��R'��F&��	�@��8�P�'H��E��KX��G"rr�[ZHK�G)�c6R2���=n:�HU�@6��{Q�f�aAb���<��װY�O�}Q6�w*���3��#�����I?I�f��>�%&>4��y� ���VrCｰZe�|x���'Wj��i�o8��e���V��2h}���=�)O�Qe�F2�!�45�L�4ՖuVj�a쫓ρ��j�+$���L�����BU�{�^���T�� :��vYI���
-str�gv�B{t,����kk3�hƃ/�I�'�_%߿��j�v�M 3�ѓOM��D�%�͸N�������z�MD��+���z�@�wL�5t2��_~�c�E�7��G>�w'*3\5�kImt��m���~Oq(^�˘��W¤�z��%7���C;�j����p���v��^N7	a�cz��u�o�j���'a�$��%�7����fQE	6c�c��|Π��|��&� LD\������Pu53asE���z�[_�&�W�@i��D�%���Q��kA�_�4m\��T E��3:���ÄGZ	�@E�YdF���-��>?s�Iz��b��m8�#C[�-�{�뢢!t��!���R����g�1�z��E\���Qly��1sF�;/
l2��g�(e����2`�����H�Bl/!� ��ޏ��ǘ����M�c,W�|��8d0+vP�]$B�v"��GO�����+E�a&$���ћ�P:�>K�P2kŖj��0ߘi������L��o��4�Y{y^t�<6:�V��\�{�}9I~@`��;5�W���o���j�9�ѩ�Q��t���]���k��ΐ�M�7�D�_8�<�C%�[<2��� q�J��ڂ'�B&܅1{�h�����pg�-�^�Z�����*bA�ʭ
#>���+��Bn��d�bksx��x�#}\֜q����|m~�:��'U���A�V-���8=�P*���]	��Є{��9p��Ɵ\�m�ی����o����|{x�[�h����k:�h�f6�>߂����j����<�'�(k�p4��V�I+�$���L��K�5ʿ	��J��l4���t:e��<�9�PU6D\�j��m?[nNp��)�7��.��쑙Q ��uA0��H�Lm��P�ݰ`�1�ixʧS���\a�Y� �~����i����.������|�ɜ��V� �tJvLv=rq�EZ�0+�R�b�nE�G��S+o�V��)-��жx'W~�>3�_[�x�����}�}�z~�ʃ�cQ�C¤��-	 �"$��"��5h���K����g�k�e�$Cjk*�XE}�>�~����וVBVk��'UR>�S����r6����8u3�p���FM}�ԟd���d�n�m?vR�ܼ;�?�~!�l�9�������Ti$�	�vp�}�����>�CөP`�^��,��]�&=5h~�O�{G�O����[�$�G�r������:7Rv�����IF^���9%�L�;���l���&�z�0,�Y��-S:�$���f�	9�)X����8_������O����9�O�k�塩\S�m���B�+X�9�ylI0k�����C�1{�^�� ���-4�8[��8�5N���I^J6sA����ʦ����j�QY������硖�k���M�(���_/uu$#]@�>�$�!�!����Ea��=����fw�>H3�94�Q�]!g3v6*݊4������ǥ)����t��T�_�P���6��~�a.���7",�U�K:�|/���βڶ��]�y�}*�?P��*�~_1�y�.�<���%�L=�-���X���>Ҷ��*M=9��P��od����ck%��x}�ȒMP�I�]	��1mS5�Ҧڝ5O�`L�@卬F�
�%�����7+Pۣk��I��,�G{4BI�0�1�֍�.�K��~��h0�4�E���;˺�~�{����,S�Ѵ��i��=���.%��o�˹�A 6��Z펩��Í�ݿ[�q���9�$M��<q侺ň�����+���������=ʐz~Ffu�X�|�?��}o��K�!p0���ur���8�lD��g�T�>�P7�����a�"3d�3{�
g�������J��%�����|�_#��N������f�j�TO��9=+qT�6�#�L��vf?Rk��|��g���qm������O{�֦<���K�ڝ�E������(u��տd�!�ӗ�A�vi�d݇����f���i7��тG��C���eCX0�h݀��A����'^X����'\�eP+�θz��J��A7�K� u����S~�Z4)��p�W6 �����$�+p�c����`&X��8Q�p��w����Ϸ䠊9�6���A�H�ӗ�u�pV���*}���F���x'�ssd�����1c���{�L�z��R"��o?E}pA����򩓲��Cʜ7���*G_���cv��U%[:٣����|��&��y�|����C�w��fv~]��__�F7H0���$��p<^$��E[BM8�NEG^&�ht.�C$�Q���l�uo�޺��`�4iM�w�q�j���cN9w�5u<ǹd'Y:��n�����.�m~�}S�֥���������x5S�-K��y�����5]G�_�R�-��x`P�8�v�(O�>�n�ݣ,T�XQ����w��������� yR"Y�#l5��`_��ݍغ�G!��f߅�jV��+�����ƴЅ�����
����=��޸ �*
Rj:m�z��>�XS���=:��uy��}F (@�ɽ �X}���p�&Ϩ-��a~'��J�'�:�\}NP�U�&ֽ�m6�n9B�����Z��+�V�[�=���:&���H����ʄ����wR--VX'����kT�g/S��*9 ��T�x�r�L�����J����#v�j15l��H��`����07��gQ-!���@}U��#ƽdL�6Ά��
Ȇ5��?�k�2C�r\`q՗]��b�w���t���yb�h�&`�!�+��k0x�í�ϛ���J�{[K�x�(u�J�Q���j�8q��j��@]"���z�8e�i!�#�Y�Y�1[C�u(��| WuFR��}�S�-�ƹ�0���Q���.�6wm[w$��Z��C7FMЙ���o���ZTnSfv�-a��i\7�φ��_�v��i�u,�eV�;�'ᶔ��B�	��s�a��5g����'|����%���2��\1v�Xk��_G��!��a��H�`����*�41`�~�u���cɈ��t<�	�b����a���0�$��e'1ί���e��c���
���fjg�*�c-z���m���ٚ�����a�fV��ߏ埞�7��-�cfN ���ˊ
��C�+��a��Ѧ��#���a:=i���ݦ]�W�ú�{K6����*�%��d���.�7�y3����-�ʸ����G*��N�Ѳ^�����}L�[��
H�9e���"#Z<��
�F9�6�T�B�ix��P�_�3�̪���W�f1[(��O�|�S����|=�$���b��X��٠�f���:{��J�p��j~��,��-ST�z
=C���+��}�?����X��-�H�k�~�}��XD:I��
�q�h��Dj9�+#D��Z83��På��{��K�?@݂�uq���Tȟ<���J9�!l��|�3#́T�T N_����"�4?���i������0���`����1�n�=�����r�(j�!H^�wp�e�<���\����haBxPXFiY%�Sgd�����f�*�ZH��ɩ2����tƩ�*�(RU+q�h��z��h��/�)ݳ�P�c�SPs�H6���i31�~42�x�Of��l\,���\���x}Y��>9=q�ґS��U�.����<jK�l���l1�#�������m̲�����X��u��Ē�)'�Y��G��}�e�����ū�b�3���n��o�\�G�wį�/m^��P0n�ө\��r�(/~�=4,��.�姚�LCn7AHB�٫~�#�y��cl�qt�*����ApCZS��.fe�s�6������{��BO�<ae:6텖S��:��N��.�Z:0�ͣ������o�(O�����'��f�y"��8���M��q�U�<X�^���>�!R��q��<������z�V�2"���s0�_�5E�HJ��ʿ���P�,5O�!��1��X��7Fq��̔$��j3��w� ���k��[
7��<�E�Ӣ��~��x�B
j�y�I�.yIl��}�-ɌNR�?�$�
�����&LC�DfP��R��J���݆�׈O���Ά��/���,[k�R�yEaQ����3[Ҕ�ڪ�B�l%n�k���@�K��fT�
��ٗ5G,H�ߴ�6r4�id�LB�O�[�j.��e>��f{ġ���@�Ñ$����'���䱳�yl�sZY5��s���5����k���7{� �c�Dqn�C'�q���Љ��S+)1�I&�4W����+u�8D���w�ʴ�s4�Dse���;tQω�{!H��$�����n��P\��n�y�m?���Z.�
5���%���+������/�"Q����K�K';�0+�O_���fpm�ֶ蚾C[%X�Fǳ�	��k��p��/ 5���Ge�K�;\�R�+��2)Ʌb�S��&�kS��R��%>Y�'�M������"��gֲ�����j,���<�K�p���Lz?���(�h���p��X���[zeON��B���J���qSZ%�;/SSr�A��RO�>�g%*V�9K!�����,�M���F�� �ね���ѱ০8��r��wa��'g'���km����G\�Z�Y3:��#�Mp��I��)V�f�֨���ˏ6�z�<#Y+�3�=Z U��Wں��-2⺃��>Ur��|֩^n��n'�Io��D%	Nvr���f2᪣�L�!JÞ���7����[����̖�����SL��tGy��i~�Et��TB6��O�Bz�-V*�A��o�Nb#W��J�,�W;�EZ�h�~-��:��
�H9��i|�
��󝾶Lw(a�x��ZG�(.��<� _�;dּ�5<�?C6���[�D~p��ep"P���4\a<�|�E4��CLT�Gz���P����6~)5�^R��4+�{Oc�m!��U@��s��~#���Ygw�Q:{ԄDA�Hǔj��`�l���m�z�T���^������(��y��yo9(^<iJؠ�X�D�H��~3{�Ze�hz�A/��ܬ&�L� �q�} �#j���U�ea����m�~c��J���l�
�R��3U{��a@ej������7��U����~kz�j���vi��&�h胃F��%=��o�ETYB��&F��l.<?�-I3�t�'aV�D�^�$�~ř����闧U�p�$�d}!q>ah�Ă��~t0�jn����#��)��Uqs���B�����	RH�	Z [��������U�;Lq�t#�*��9�#gCp�mX�B��bj�U4��ݏgY��,�}PZ+���OZ�YMh�l�dH���c1�]�tP-����
�jQ JAq8��|��Ҡzc�Gh#��p|����2�b���QI��H���;
W����	[�e���ALK-є��|�L8Aqrp��s岎z�B��5�Q��0�b·��5�X�H��w�~f� �i�p�Y�~�.ஊEH�4�/}�J�hu�[��1��k/o��|�ߊ�d�cf�AcpWq�M��oJJH���t~u(]�ݚ��F:VV����GL����4��f��'�������G(=Wa��?��)7���`{��P��s5b@ɠ�4	�03��+�߁�pߔWH��^�M%A$^9�>�L�o�NEt8A+�=�?1M�}a���V����ϥ���l�'@a�dI#����h!�H?�M�i��Y��Q�m�y��Sx�%պߙ�!�G��0m���ɓ(�B�n:#	ڹG��$γ q+�x�Ɋ[dO
�)�@y�>yS�-8.:�=�W4�k>�f&NWtO`�^�57H6f25E���vi��4���W��Th��� ���eۣ�ub��h��U�7V�7j��kc�{u��M^Ou����p��}�S�t��KSf�`+�5K�F0��G�-��ݴ%q����2�P��I�D�����-��?�i�j��"�lqln/aQr��[���]�d�XL�B�O�H�F��ڽ�ϣI~�<�H�8�q�9w����-pcRފo�5W�����6����y�_������yhiu/�pS�(WQ!�O��hn�@���r�|�U�Vfٛ��!�㵪�R�+_���6E�f"8�i�)bR�w�p��X�rҹ4�؋�t�vDU}����ΆCo��#���X:#9�.�%��7!��W�d�q�Y�5v[&!�/6�a���&�}Me���5��\�a�$�K3�=�Z��K�y|	�x)v��3h
I�k�8[���CY�9�"-��b��ʲ�8�!�[�ed�Ρ?[��m�gAX��Q_2!�2]+�*�^���_61��ΐ����F���c]׽�J0��;ad��n��|43X�����?g�/r��h�?I�tf���X�f��N7�i���:4�շ���T9�Tɝ�l	�%��5�J�@ա2Yg�t�<ԕL��KO��W��|І"Q��[97�b�;V��K��F�]���}9~��-�
E�AЅ8���e`���5�K�5T�-�J
�� ]��wE���d'�X��Y�{L�Ͻ�/��pd��Х7��ofM�$��n7�n��ƒ�P���z���6kjMx�>!�O��G����D�����do�� �����}v�zﺩᩋ	���=�05s�T8��x���T%`������f�P�F���1���i%�˥�9�`\�&�����Y�s����S�l���k�t�����|rZ����$7���"���C ��	�]ωs+5Nf����0�?t�k:�V�@j5��泥������hƄ��m�"ywc������N+�wa�,��6�9c�%��J�Q ��qx�e	�;x5��������HB�	���$��#*����v�յ�?9"M(��DV~��Z������N�^|�k�S�B���Ch�0�'�	����ŕn�dc|��`@����=���p�NkWm���F+ox�l���@����U=�}�Q�7�I<�`2��� ΑI�R�e���L�J���gA�^��-�ˆ4n��O)@Y.���߹�*���?nnl.���,?w{�e9xn�c�#�g2!�����ԇ�p����� ���֊g�n6jg�ݤ�D��w�k����<B�n�w��ۣb�=��K����O^X���+�.�L͗SOYf�j) �"(�����3��_����L>t��aݭ@����_��X��?�Vv��Y� �\r�B=��u��7+_a�\6�Z����oy�{߫��I�r�����{�<��	A^h�ha��,9Nλ�U��̳����m��fx�^].�`kq�{��y�{6��	���4�!��`��nيSe剧� ����|ꩧ�� ��yh����Zy��U�c2���7�?�,Y�D�z��������؈�E���}W�k��rQ�Ni�\���0����faiٿ�[3xӞm<W����v�1Md�̦$b��6Ԧ @������ܢ{d��sn��`�{3���fdS���s�|<�	�,���eB���mA�&)�x.6*aͨh�����Z���7�n	c
@םq��N*��e��?��I������#��r���m��B%��B���=�a^LJ�l �!����ݽ]
���B\�L�=���fM��j�a�[&˫/�B^{����PA��)�����G��C�ۨO��c��>�6���+L�I'��e���Ym���������a޹���y�0  pL&�(�ʠ0���c��]��ʕ��l�/Z�$�d���+�/��dD.�u{�r��%=��q�O��g�cNF���C悈�2��m���0.S�k�<��s+M�j���)`�`�N2V�"�9Y�Ƶ&Ș]0�7������6�8�E�(x�
�;��m��� �� �XS������/lIg��m���e}gW�(J-f�H�`�H�b��@�iZZ͝�/�5����>�Y�H�U�fLozӛ�G?����|\(8�:H��A�� 
a�1΁�q����{�9���uP�9|ͱ�&n3�!���VѶp,�t��Y|��CK�a����I���h#�YP+�y�+����ʍ���ovъ7�&Յp�={�Q�^�8�S
}�R�`q[�V[�y� �nb�?@��o���<�DW�[锉u��D+�� �mj�Ԩ)Ad�\ 2K�K!�j�Ԩ�ٓ�������S��B���jx>�R�pKoP����s][n����砐!S���r��D%��Z&ǘc;�)hf'�E%�S�;+0"���9���)Ӎ��Sk9�N)�ӎ[_c>3 �$��U�Vi�}��>4z0v|��|@���AK��xZ�ZV¬'Xp��M$��Z����Wf�c�!4�
���`�3�`��orB���I� C kD��=��D�Z]0�0AH�:��4%E��9��&S���q�>���Ae��4Z�ʲ����{��[�Fv��l62�X�ڪڭ��S��؅3�5�	�^1�`Xd�7k��[���1���9q���q�ݾ
��ϸ �}n�}U�c���?X}�|l`ι+�"�u�jSxP萑��\�����cxM*9n\�֔ƋB�D���*�V�}�>G���(u��.>$UyAY3߳f��x�L��@�(iM�V�y��k���Jv��M��.�}�z�ɚ�w/��:a�����^˶`�c}2>B%�c��H�A�������<hR�YK���Cca�F���# Ԣ�_e ��&:M^jVdH�	]F�����'�9�	�&7L=������L�Z�ٔ�4�8���2y��j,�}{wjuC<������c�\Ư��76��zfI�C�ɝ��(�x97�;6���q��Ժ����2p������$L�q��]?�мO��.�A���i�3��j�T�sq� 7��bl���3�q�C����z�TɨR0x��n@V�&ok����3g��!FѪX�3\: d�gRz���ף��F�fQ	����Ý��|Í�p쨔a����G`n�t���o� �7T.�4ak���ΑF��e5@�'��H0X,$�KޠT.EL<ה�����ӛYtA�ܰ*� � ��P�Z�|h2�Ajl�ri�R��Ak��1Q�@��}�?]#��
�4�kt��*8��s5�cw�i����� ������OF�Vo�68:��}��Q%V��;wFnBׂ��B�G�w�n �V�{b����.��2=� \�َ߃\��gD	�p=h�(3 !F��Z0xKbk� �lT�G�؏�DH2/�����*3�Y�ZdAֱ�����ڗ��S�k�PR%ݳRƒ���c�*@��芳�����z�5:�pc�0���G,�`����	�*�q�tsj6oh�R����M�h��z47DD��0Ml�FZ�į� D���8��R��@.�!���q=�H͎.�Lʞ��&C��v,۰)ߨ\�ճ�`��i��/2�t�X&<����oW�4炕S]�>��=�c7�t�n>7�]����;2N0�~UPD���
��Z�h�1F�}�_q����~��������8'��abS��x�-��d<\fH0��,@�0���	����������߯y�k���>C�_���� � 0@�l��Z/A��6��BU�޾^�_ 6
����V��,4�?~��(yYM��֏����
E9w��7ܠ�?ʺCQ���
~���댖�Zfx��s�X��`L`���q�����f��v����L��f
_A��R��B��G퐈�������Zh��k�>{����]��ɧVK�*}���Z�@�YlQ�ޫ�G�;�O"+-��.4-)��) Z�T@W��v�8�Mr�>��`=@��&eB	���q�\��K�.�x7(��+�g���!M����`�{隵�ۼy�BfP���KK��up,�{�'��\ (`�x�5e�b��!��KZT�:��"����F��{����u��S�į�_��g�2�W���rkn�"�g̷E���ݣgq������ *JVٲ�����B�yC)g�E8�T�xp��+�d�a׭��v��B��1*M �����#�礹Z�;q 2w�(�M��Z��+�B�ߥ~!��ν��COjUO�=��%��G�n]���f�$5Ϗ�:�7k�'�#�%������_Z�{��H����6͋[eQk����܋-��$޿�����w߭��:9������&����`ʌS0���Ƞ/��zX8�t� ��f�ƅ@n^������,�×���~���Gq,�����gsv��p<~ñ� �|�I٢�O3v��B��(@�U�u��SOJ�-Z�y��ǩ+4O�e�&��0 o�O����[��`�"7�H�����q�� ���`��S
�M�Av5|��r%u܅� #�@�Ƥ�ZRm��=��<���mL�Nm6�|����n��֐�^2�-���������� ���F�]�IYa��H.0B��B7m,%-�e6=��BW@b79j-6�4��z}�[%�;4�@�k~������� � ���C�	\�0?���� ���r���eP��Q?� 7�k�cG��!�tAo��袱L�U��k|�\U$��2o�+�j�{�N�/�F���	_���%t�Kk	h�����0��ZP�h�q�k�`b"������Bak��?��gRҹq!3�B���es��@n"�L��Ԉ�v�b��ohz����ק@�����\��B���6��w�N��]Q]=V`�B�n����_ށcC��9� ���h���
 �#H���g~�_����0��`&8�����Dt��."ąC2�ߏ�i�L}7�׍Q�� ��pqshE0Ǆ�D�ؖ��h}�0O�/QP�s��5�ǔn�1�u(��^`��5Np�:N��3Q �|}�b�� ǂ�(c@&<��ts<��606��/Aᅟ���TF9wno�C�	����΀�3qӻAN,.|�=>mdsp��:l���.�:V����W얖f�,GG��� �y
}eim�&۷�UV�Ug��:�4�7�X&b�� �(�_{0&OA@���,��l���Q�%��5]j�86;|��3�b��,>�8�b�q-�tuv�0b�<|��l:Zp���5>��I���q< ��d�8����?�=��83�)p4���\�ŭT�ZXcO������9{Y�v=���B9�bE]�%-����C�K_��&��Q����z�9@�C_|����q��P�y�_��7���+����omrq� 6}�4��F.$���k��(���M��f����Ѓ!U�[�R�5&j�4�=X2]ʅ�m�e���Z�X��*�Mii$��w!c���3�ʶ�.���w�[�����I.y�7F�}��`�6���\p��Ua�a��
��[�S&������`� O?1�y�d�T�������k}�k�q�x@�L���7D���Xo�jH� ��J�lI��1
$�V��gl �#Z�`�e,�*af}oݺMv��"�]����݃]M�R���e
J�) "���泮C?���T{���\��J�Pֿ���u��O�r����:��?����#C���T~�\<.' ���+������E�z(��ڵO�=��J��\�Y�[���
T�D�K��֠�. ]L��,uiycMsHd��w�� ���|�)2�?h���oFv	�
����;������#D�v�✘&�����*�87�F���:��lὕ����c�7�	��V!MW_}�Z@���q#c���z�*���O�T�&ċ�̃���@ny�������2�I������c��@c?[��{�V�\�x�\|�%�kj�b����Ui��|�H�P�����B?U�NGx���=��c*�+7��E�h���Z�J���*���\S-����~�'���#��-�j���6Lm�I\<�\��bc�*	Q��N^5��Æ-Is>-My�8У�/� �V�`���m���O���>�}AK��A�:܅ձ����/��PD;L���,Y�9���
,;�5`l4�/���'�|R��c�6���~����y�E�
w\��eR�V���$��K$O�m�����b��\Q��н�w�Cq�����d\L�" =�� �YXXn�9 ��3�0��k����.����|�[���Q������/̾��%G��_)�TE B�GU�T�E:���}�,Eb�=,��P{8�󬲩��la78�Y��M֢�2���������9V˼c�����C<(�^\�%f��N�+t(�2���ɠ���'/��n��C#hmn��^q��^li�k�n)4o�0P<�}�4����Ȏ۴�+�}%�fWC<��(��ۆ�]�2e_q^%b$�p���!�l�fq��$����+��@Ҿ�V�,i�(�b�����j�Ę��4��e�Wv#J�>�'Y� D_4QR`~``�`R[��8n�����׍��w6�p0OM�:��A��q5z� 6e.�U�,m����_�B	��Gg6�j6o�$�=�Z�Ο#���&2}�4Y�dQ�L?%��T��L�h j瀝~�{ߋ~�~�!��@/������#Z�T\p�w����)p\���I^6cW������^�sF;���(H���=��@Qjn�*�Y.��1�A����\�W��@AT ��c2�xr�)��+�kk�Ұ.1��vݻX3hԂns���u���e,�>���eR��C�\�Z]WPf�e3[m�\J�+��P�y�3���>ʲk�G��k��FN;����rQ��:tĚ>}�E\��`B_w�uZ��6�x �IiYpBt�d�1���k}�|��u1V�}�g2ZO�%b�� #�����;8��e��k��$�*d� l2�M��%�nj�����K�:JD��&r���w,Ǎ�!��H����(p�(�+������[*J�P��x�jts@ns<#��<�PD����V	�נ["���-�� ���};d�]j�s6�f	޳��y�	ZP�J���E(8� %��#d�z��}l)��ZO�ׁ9����#����R���׀򁜌׾�r��F��۩ �fË�v���5�'g�q��6�w���$�,��Ϳ.��g��d�Ye��^q��r���F[��"۷o���{��Ӻ�ʁv�9��Ur��ʹ|����>�#��b�]�9>Wl�!�/#ӧ��Ν�d���֔kֆ�U�Zj)ؚ'E���i2�Qb�fj�����H��"p\+����S�fi����X\+�����x��P
���j��j����V���g���XC
V5o֕"���	"���ȃ+}��``��`~Gȧk}��4�9V����B��92T�tQ�X�:��/L�4n乂����VY|�rm�R�x�W�\�I���S5��dI7K���h������_��_���B����&�ʤߞ�EZiHXl��񤣳W�|�qy�чuMa.Qtn���SVi>;���<���Rr�D�b��{�?���̀	[�p��y�*-�Ma��r�}��R� K�_�Z@�`�c`����m�������vO �#,5Lm�f=�7����yg�M2w�B�>m���K��κ��ul]r��À�ϩ�9�?�I�]�>lb�3w�2a$��Dl����1��A7���k-���R��V?��ƅ��!_C��HVz�pu\���� �u�� (�6N�r7�}���h�=��w�c=:�>6n�[9�*���g�]��D�j��=e��*֌��ڦʱ�N5V�d����J;kR�γ��E���S�yGa@X���1�p��1c��-�o�p1G�c��Ռ���J�7��=&;w�0����m�7���O?a��.9�3����SČ`Yt�t`�;���h[�dB��x�J�	�	�g�9�x꼱
:�&�+�}�fО1��+{�w�r�u��	?�St1���2W�[���Ѩ��|�fvw�����d��=�չG{���,r4}�ثha�r��c��m�c�	ƅ&:�h0����5p��D0����̰9Yր��A."��&�t3��Aӊ�@�B��tx0��	 ^�&�L
�=Ρn?Ϗ����ʡ�?�!f{��E�!KL@`�
�O�����H#h��$Jh(ˉ��D3
Z���Ǟ���}.��1��P֘@���f�L6L�j�)����K�h)���z��%��,�[�����1A�Cq<}�c�X���Y��D�pЧ7(w˾����m�Q�ɓ��W6��QZ2���+=����+.����Y�Dݍ��)�!.���'jIg뭫C�M�F�L: l�s�����)��z�̝�n&�7Z��P�����}���
�Ǥ��؄��N�5�&tr��sf1���H���0�L�f�I/V ��u� ��0=TJD�K�KA������e�����S2�K�/� ����7���������N8A��N���ʏ�# ������=�I�e�9I��C����o~3��Z|X�lr������k����w�|��%�i�����uP@Q,��}-�u���J�{�U� x=�����X�F(V+���f�K-�ַ�U_�������{J
�����Z���:�%e��������M4_~oo�TM���^������[.X,��:S�S((�z���@�Ρиg�A�HPH\�S�LW�	S)϶jKy%�:��h�6�J�5��.D�{dR�$ٵ��M���Z%69zw��t�x��~�^�E����NYֲ��im�I.m��r���E�R)!���o#��Z! �XOl6�Q�o�� >C\4�0@�.�G�+��:0Y h���+TS���������|�Ҙ6�]���2�pʤ�
�۷�h�}e�+�����w�B����5�gd)
�qpO`T \�)��������5F�s�O�	0B������
��A�J����j��]pġ���d�_��v�/�˥�2o�!�cm��P4?�s`�̜�D�F�+�i�T���s���SU�?.�7˖/���g�8m�Ƿ��-:�_��Wt�1Gl��?�vwȚ'�ŋ�Ȭ��e�_�4���^�3�=�roi��Ï<(�/]a�grdMn޼�Go�3͢��2P��ф3ƎZ��93�6��l�~�L�fi�e5��VnՒE�Ф#���7��C��\D�?�zܐk-mi���'�o�M�ךg(X �{��- �?c�\'1���h7!���nA5$>Aಅ#}���c������������$8�52W\��MX�((x#@��+��2�� 0Pi��#-���&����wn� �k��q����_/pK��ѳ�>��G�"�@�k%!��6r��D:�@J"�@a�u���%+��_���eS����e��Ge�	�$�d�~�(�j�%~�C!¼3~��}׮
���AX������K��	�פ�:��;�aƻ��ת������̄�
%��n6s>$
�:�q0~�q��=p��A�ɕ�If�E��[�[��,��#BX��Q}���m��_�����;�!g��)���m�ҴԴ�=#T����O�T4,�(�,��%}蔟Ua�����C��J��)*:�p(n������}6wN�4vb��2x���، ��]�	�bW��0��i��������<t���w��C����Ѳ�𾨀pL�}���;��#�{�6D.�����8�pq���RPQ���g�\7���<����p2T#�3�M�6���}u�jv���X�3��N�9k��q����[Rf���=���c�v��U]�{h��Gy$Z[ �0���]�7�e�+����	q,V�| N��b��?�y]������Z�{���}��0���o1������f5�b��S9�M[,9
Be��S�<����� �!͙��f�h�A�*�XHnh
�|.�Bɨܶm՘�״��V|iknU���#!�h��Y��|S����3���G�K%V�g�?d.�r|>��*�4�[4�-pr5f�,1=O&��{@.�хK�̏�w�%�(-���Hp��ܠ,����0��ɀ�c�2l�QQ�x�i�1�D.ѺaN��=����C#�K����@ �4N�ux2Z�1�^��a�a_@1*h�W6g��t^�����+�j6����X`�yͫ��y��A���,�����
���w��	�
����
�2u�qъ�eZ�Q���Y�ip9�I+��9s��!<�2�u�憛��?1��PD7 &�����6���=Ř�U��U4@5%��)��}$PuHW_��Ɛ��877]�(I�m5�!x-$
�ǲ�O|���1Y��t����b�5�͒�޽)�z�t#Д�2�`���M.�����9�x�.��ޣ�&q3MyW�e��������Em��Bf��� *�-��
>gv���;&�1a�P@���ǭ��<�D����/>���?W耈v"S#�g���
5�1�C94���*a�J���߾T��7J��Հn�Q�̝ky�����29mʲn��޿�Eo�EF!	�f�z���h�Y�e]��.C�M�k>���=�ܣ�/�ti	`<�Z'ˌYs/i��gsm��t�î����Im�F �x��3T �,��6�����z��?���v����}{�q�d�tvwȹ�](k_xFt���KS�h�d]f�m�$9jANҹ=2g^��d��ps�Իꪫ���D �����N����(&p<nb��&�M�����}��K�Lj��+����V/�@$bf����"�m�X�~4�u�nj�.4�ڸ���.��L.�P]+­�J���&�1^� �fܺ��5;W��o���� �����(���$өU7&�rqc�u9NC) |>�y\F��	��0Ǆ��Ұc^��B���R���9�|Æ��q`�с���d��^[�Y��ß� �$�L�9��0!�hˈ��4)�w�F�v�ؿ���kUY�AY�9>�' �~��� . ���K˖� [�m��[v(P��y��PpSk��O�5O����j��=,��>'�]���R��~0A�>���<����<��cr��UƼ�&}=�̝�H6o�&���/�*2�\�Yc�Z�ȢE��Y�\����{�N,��/~13�.��ԟl
bLH���vh@��~.:5+添d�ֵB�O�u�����tQ�j!�]MS���tv�� ���ʨ�[��M�'s��7�C�k���A.f�ǻ�DfF�h�E�Z_�8�v���d�|>���j����
@WP��Mܪ�'�I���q��߱E�`;�]��q�R�G�%�g�[!�E*���3{��s�z��^:s)�?��ޒ���<u�t	�e��
��ɀ��Lׅ�Ak,��)Dρ����>��ʧ>�)��~����H�s݊ p}�֚�|�lE�tv�ɶ[e���77	�VI{n4�Q���'���3t��ث(���r��R��_S�!.@�M�[o�뮽Fʥ@��Y �k!V�?��J\$U͘1K��XN9m�6�����[�zu���O�G`����Gsh	`��>�� ��!& �VS{��r�@�y���ӹ_U�\�G�v�����d�
4��2|�h�hM��ۀd0��.�k� 2
��e$W@���x\���s�)��!ƙ5\
W�P�PP��w@�_�}��u�D�w�X^�.)

�q�;D(�-�x�P�k��;}���U���:�@72�0g�8��W(<𗷷O�Y��j= �����E�Sr�+��+�`&�X3��в6Ϭ�q##w��._�ׯ�1�5�\�l߾�X�}�}��������z�{߫�$���]:�)|���_����2c�\��.Es�<����#΀�����rs_S���+*��*R�DP=���o�3���!�U=Sv�L
�&!C���.��~_xѥ�?{oe�Y��>{�]c�IwzHw愐�aPX��̹�8� 
.��\NG�\t)2xQ��W�H!!�$9@�H��t:���w՞��{����U{铳���*յ�7��3��ɮ|���A��� ��l� )����[�����1 �!���x��b��w��k<��M7ڵ�^�X �!�.��m=��-��up�+;�R8;&���%l��Ш�w�;x���-��m�52���aOeSfIZ
�Єc�^�ȩ�6ŋELD�DL�	��]�G�2AYeo��@�*u�T���!b�F���k��*Z�&5�Q(c��)s���i�e3�B*u����F��Ԥ��9�R��Ɲ2���'ռRf�k�~r-��2?�f������v�s.�|;c^Fs��9J���9i:�j��y^��C���G��7�ךA��מ�y%�s�yf���J��9��V��V�c繶�����x��h1oذ��M@�*A��_� ��mp�$�~�sx��\?�?kn\)U\�'������>�r���V�6�\u��$�YPD�	A�B���W9ae�4�O|�U��^�:_L�߳I�� K��ˎ��O�Uw�Z �� ���čMQ
l F�{[>��NMuY�)m����("�
����~"��k��Y���MoT-�)������W�kP�y�G��|�jhb\O��y��R�M~�7�c=T25Ʋod��
�@(�c(�bl<���I���¡�Oe`�!a� �&��0~1.�Ȼ� �^x��)�)�nP�}�	s���'1<1/�m�w+�5�)H4_�#�d
�;��(_�y!g��@���wx��pN�A�λ��]av�����	�2�hS��iw	x+���,�76�s�O�B��u��(M�g�p?4a!H�W\�_G��6m,۶�[�λ��3�mb���pѿ���v�|�8�,*��}���
��b��O�?����ߞv�Ev�3��o���i �$p#M�N>S�3bʂy����ӟ��8t�v���O��o��661ލ��s�p]\���z�T�{eh�U���n��׵��J��C����an1��.�A��.˒b=E�������!'B������pec���k^�':hD����P�5�%�=ER .��'�t!|��_��\�/|�δ�u�J =/{@8�t nDm8��Ĉ�׿�-�})���H��`116���B.?)�?��Ow�������b����"��\!"������'?��o}kW�L5+�M���LEH2�d^ٷ�SjӀ��¼0.��QB}���|����Ks�&��<�&�Q�{�~{��;7�fZQvdHs^g���N��K�p�g'�F)H�Յ�Y8#�S ��d����ǆ�ne��h�n �L��?�|�㡞�x�A0_���&��0¼G���ёh����u_�[o��g�$ʜt-�������������:D��<�h�>_Z������i�س�������wo���ZR�zh���V�~a�F��DȦ�T��ɒ��*t�<]h�v�i�>j{�;<;�\` ��o6�G��=�K��@t�Z��7�Ϋ^�*�w���*�A�%*VyOȑ�F�Ď�Di�H&���qe�� e��3�xS���D8D���!��nਬixaF)E�*ڗ{!���Y�� �C��<�@�#y����(�����B��W�W6\){?�a0A$<${"��#80؊~���=E�A�T?��O�{��^+^bh4�94	4��%�u����&�>�\�T��h�t\C�*����&AP&�ά�C�e>髊�@�`����s��΀�?5d����<}�ޙ[�瓋i�����?������v�3.�y��.4�hƌ���Z��f�_tG�۲�ϱw؇w�xR>��}�s͓���P�%�{�� �� ��D���N�CoP��Nx���uVe��$jB5�i^uhI�i����\��o~�C�!<"F��H�z���F�պ�a(�i���6?;e����>RN�P�s��	�-d?�������AܐH���7T#��T`	6>Ă�90�*ϒ������U$Z�	� ����1�)�"���4���B��Y9�"�����
Q�@s?��ϐ�d���B��{�~q�G?�Qυ�Drg��P�����{��!�H��)��!
��9��ClIj�X�]���ų��r�i�ar�9a�`�h*F������u��z��_�-	��2Ϭ�`42�0P�
q���_�����m�Ͽ��?��cR��kVwn"X�f��:�<�X�AVd��\J�� �V�y�~T���ce]�3�XWi�eQ�W='�j4f՛��꙱9���A��d�	O�����R��O\������K��n�9�HNJ6
B�懀�i{SW����������o8����ol
�8
�d8\��9x�"�mi�����7�CL!(%>��!=��#M�BAuVrۈ(wp/s1�:$q"D)�5�ZE�
��D��k<�k���@���* v܏���X_K���a�1	P�;c�Y8@�t�y/����ғ�E�Y5�-�*/2��nC�@�PY2�DK���Nt��%��w40�>c�Bg.y'��0�Y��~�E�+h|��4h^�	L����ݚ=�c i�B��ǟ9r��*�! a���:�C�AY�琺^�h1�s��w��?�A"~�7~�mx0`L��%�F�)�UB{\�����#f����M��'��N�6��I���I�"�r��>O��xD"/I���&U�������~[D�JQ�,�!�mE��J�ǉ|!@v�j���SL�u�!v"�����|�c�C���5%oh�$�8�X�9��Op,��1�*��sH�Ż ���x����,�i]Fb�R5�hD����^������@Ӑ�esк�/��E����|(�KP!��Ar�鏘&���i��^�W~Z�]9�i���
�VQxDI�k��\�c�b��aj�����p=�DJ��h�p%�;��jt��Ԗ��,��)���t"��V7�R��4Qf[*G!�!g�����<���c�a�s�s����5ߩ`#�I��ƽ���L����	O�����_�Q��æ����}`%?�^UL���>Tw�y��*؛^����R沴EO��/mz�p���ik�w\+��7iK����6�s!����Hlh2��2x'x4� |b��$m��8��Gʂ�+H�Z{f��:�`���,-�#y��� ��Wy�@�U�F�T9�0�a�r�4��B�=�R3�m��N0U�15*s/����+*M��҄�H�Q0ϡ��1m��	舾2F�B"%��&,�Q��#/zFz�41d���\l'$G+I]P%�����t�]�fUA`��|م1�O깕/�܈KQ�V�a�SGm<�{ͺӲ~������u�7��.ɽ���ޑ&�%��`��~�<	�Cc�ӂ>��M	�FZ�[�Q*,�?�'in������{��S�L�Üb��Z�Z�Y����\�����,I��z��m��Al�&g�!�gO��A=B�a��*C��(�=i��w|b�_ �0v�[��C��MQ��H�u!L�7��	B
T!�q��v �0R����4 ��3�:����-oY��h��5���g]B�W����p�.A��	��W�
�]�H� <����?�o��R!-b�3`���	�]f��[����L���O^6��Qqi�3��G�G�W��H?�%#��ɟ�I�����Ea_�y@;0,���3704�R�I�)�6k�=r�H�����^���ʠ�}W�����ϼ}�|�~L$K���=�ަɧ�v�yOw?�b88D�+�]f��	wj�s�6��g�䉖2�4��v�g_�m��i�^z���lP;y�}D��AF�?����L���I�-�0�I���I��,����{�����'�r!��C9�9\(���������S���6���0xB�t�E�$�*��?R5s�����+�} �G��!�Ҡ$#��H	�4���:4�s���Ic]�w�����>C����T�{�L��ES��N����n�U�A|r[Mm!*��� "#kߤ�f��@' 1�h�N{ы^�D��q��I��Aȶ³���=�D�1��Þ�d�D+�ko��-��&��{���	�j�����[��@`Ew���<����&�sS���]�ў}��8\p[Y{�,Ac���pX���h�Ae<���$�)�Ms/�w}���|�z�t&����N�2��Z�W&�7"��7������2���#�
j���1K*����q�/����>w�ҍ���f�o����򐧞&�9��呲5���a��ݞ�-�Qbu��d�4����aʁ���W�b+�'��0�Bd��!���NW�p�ͼc V&�:��Ƚ�T���+!�+	i2��M�7i6��& �5/{ُ{��/�K����9��D"f�䨨bދwRn����e<���K;����L���@��y�ޘc4i�t�w7�|��^S�"K�Y�xўpYe� ��V�P�n�&��Ǳ��C��N6��7�4�3� zu(��EQ�S�KEzt&5\�.��pv��m��aۅ1���^j�X"-ƥr�:W4i`��#���8�,� �A�R�u(!�xSc���_�i&E�=����OїZ���Ķ���V-,8,�CN+���?0�v���61J����*����r6[mXeh�#=Z0W��!�O����$:`y~�w�c+��%ɚ�a
@H��4���"�\)8x� �@���K��O���k�%sL ���X��r��; �MP��e��zJJG��i gA�!���`H�e�8;Fd�A�af�*��@3>�x�≫!^&bN41<s�ԯ�q�T�L�H�H�w��6�w@r0!k���f�5<�5��9Zo���-�
�G�O*��N��bVr�;��/ =@¿��!��5�U��Ԑ`���eƤoT͚<r��AraU�G���i�9?7��[�5�Z$���,��&�E6&�����71��Z��KsHQ1�Ԁ�w�N��\�4��Eӄ��Uׁ�MU���׏B��Y�$�b�z0@��B��b�i���F�-�t�fl�+y5k$�����m���?$��Mws�C��P�š�<����Y��Ɔ����Dh	U�H�X�6Ұ\;S��á�� �a�PA&��5�\�/��H�&pp�Va�;��&� =�@�C�\!Ykp��q��t	؂a �cc W�p���
��3n ps�*��H����0R/'EKRO��@����(݅��T:�9H�0 4$�|��(���YW���,�3<�����K��K]�����ye�06�S��-�CVnm���eײ����92� ��w�C�D@��`E�Z���4�V�Z�l4�*�B-V�Z{7��%�C���=)�]�iHJn(�Q���b� }���L{�@/�?��̘����B#]2�I�,$?lj����	��V�d
o�A`+5A� $�B�� �Ky��c���������I/a�h0B�ɓ��Q�j�l���p!��Ea੯�a4�t�Cͼ@�8�B�P1�H�|�DL��%�mAϒ7�pr��J���c�C���5���x�,$y�m��)���˚DF��cj���H�z ��a,<�Ƹa J�3n�@�8���������9t�'�PAY^���L����B���鏌��v!��k��3֒q�n�
?�Z�y��~��{�\�ϐא�ni����\���{�%�w��J%h;���fg�:׫n�o7��ɝ�';\�nS���$Vp�tzv�Ƃ����Z���H���9̛9��ʜ#����#��,F HL�Zڀ�f�����9�Ym0�r��'�+�<j" *l���o�SŽ9Dlt&�Ŕ���i������jZ��e��C��x�V~F>��}7�a���Lu5�yK|c��#H0�?1iw����34H��`��[��uO%��AG�aH��n8�*�1f�_�-e?_�P�KJ����I�$Bļ*���QZר�[,��3��He��3�+Y�=� �\AT�tǵ��+�>�LM{G��$P�lْ��!�K��Bc~�b�\��()]j�e~蟼E$}
����?0�UQ"�0�sn4.�$� �??����ĝۋ�Z�<����-��� �չ@��묭�,���I�d`rp�f݆��ꗿ2{j_� I�!`�8��k9��R4.Bb3ќ��d�Sռ�`���{f�G�ќ�a���[{��:��I��9�I�b�J�g��CF����F��<0��a���`�fa�	 {���������\�ؖ3և�Ƽ�h����?{�f�7H��M�XS�X�-7���D|�FX�E\�R%;l»M��tjD��|�N��N��4ikj�!M4i�b���I����jj��ׄN�����r��@�"�)!@Wq	�%���(��Ɯ�A��T�L=���IS4{R(?\#_��&�K�&C�[���	�2�,ͷ�M*!��6�[g��M�[�k[��0ng���:�����nrJ��sh8F�N!�=���oe��,�FsL��/�˺p���4ڏ�'R�'�'"��aR���h\��	D�'Xyuq+����˳D���W��Ը(i^�&��Y8�dAA��K���z�-h����>6���06�,��Fk�I��(mR�4Y�]<I�������֞�&	P�H�B�V1K_O�C?MN&)[D��P����B���AjH�O�����.��#@�Z�`�(I_k/��ԅ/��Dr"�i!�t�(�X�g���'iB��S��i��ԦEK������(���X��7�nh.��Rv1}���GK���k �Sg�]����:�ߞ�����/LZ����({-_�.�HZ��3����u�x �/�F|y&���H�hz|Ƴ��F�?��/�$ոE�?|MB��v�����9i�8jRW�I_����_���S�/�ik���[�x��a��3��2�B��B��$���.�"�"_�^WO=�	R�߮�g��`v�У�n�X.��P;�G0~�ż�f����Ŋ{3t�����7�I+��+C�6t��_�Մ��`��萪�ZJ�0��'�OR���Ii),�Fh�����Z ��/%������Hת����;D�b�2슩H��~�@�WذRM�=o�j�� &�k��X;�W z)Õ�"Mn���z�W�DsǵbLi��U�?��_���q9+�<�y��(N�K6>6n��l��yf$;�����ؖh���B���~���C��Ԙ�6H�b�i�.�#��g�g�|Ye�䩛}�Q�����~d��ضc�×##�~�/<�<7��ц�GiH�l;�?zj���	����\eC��9j�>b���ȑ�~�l��9g���=�<zȞ���|�6m�h�~֕��#�2	i�+Y)e��$ &�jË��0�"�b��9�d\��6�o>p{x���i}>�w�˹�<(� ���&K�6��8��_(/!N��K������P�T�m�<�f�K���a���n
��H5�� �.Hc�Y?-I�i��R�R�MR�$i��\wS5=u�L��Ik��9�qN��pa�?f#�9���I$<��w'�@Fa>���g��51�T�*¥yW_Rƥ>�{-Ո�YZ�MPRz����ƹ��J�.���K]>�V7�g�1K�;�-����5:uZeO��Yϵ�G�λ�2�Xw���C6;��e!�;^��
�B���L-�e�i�]�����3�58�����k����s\�����l�Ęu5[�9j߹�[v��~�֎#�7�ȁ��/�/�؞qųm�:k���b/��푽�����,��k�z�&��)��6W�q�.�;�l>�4��O���A;��>.��/���E
%/�p��\�����䬽����D�MN� �]�4G���#.g���(ˮ����x(8ԑ=l�tf�ds�{��o�|�0���f��E|�>Ҵ���#�b�"Rq��FUե6O�KR��G�<�h�B�4��u��_�/Ҕ\H$(��K��Yi)Ϡ����������R9+�Mڀ$s��&�$+�O�	6⹂I$aӔb��� ���������jIpW�N�R!���|�[����J����y���H̓a[���{ ��%���>i�cr<y��E۹�L��-�Çp}��8��`�4B]C�Ƙf�u���'Б'l$���h��q.0nn�a_��ce��_��b��3�+��qx!ur�l#˷��笿��s�*��>��O�5���o�T�u�u����!܁H	a�ڴ��i�z���s׹��<W8j�I��,�^�L�">��J��2�;���Zm��mނ�����unԍ�����OHvP��E��q��4�4�Ţ��;%)�9�fg�!w5<E��sK0^1=S^Tb<o+2l����;����Ѓ�
ߖd)"L���EA�~ˀ�7.�"����~� �ȷ|�!�#C�+�I�`=1 =���q�$6�+��1>b��3�m��o^��)����>o�L����5������	�AzG���uAӃ%K�h�i��3�3�^"���=��^O�G�A�/A�<Y��|�#]�N��-�N�f?���m��u�ٵ�Lв��/"���f�Uw�}����|N��p>�v����bXp_R�nX�6��V��x}�ݻ�m۟�tr�o
WG�=���5[Hw@ �ݜ1|�(	S�n��'�	~+sd/,Ե�|�E^.!}�=ca��0E}���u�~/�⣶������)��.�E#�	��I�٧��޷z=z��SY�p��ށ��@<�ʔ �CH�^�c=nsS,Y�А�R"���W� I�J�,���u#*�\?xa�Q
!�������1����<�f5�?aZ�/V2��� ��q�He�Nޖ�] i�g{��Q��w=9y�6�=y|�M����]�S@w\�O��د��hIr��@�8q%ozӛ|O����M���<�|i����q�w�=g�����졠���]�r�ssպ>r0��z���n\>s�9�o�#�|�=Y���'��N?�f��2�r���b����8a���I� X�����{��zo
�0(=�`.:v�d�=��!'`"n2���4�}"ps-�0�`�>�'�=��s��.�;$q|�\��绑�MWg!X4�#�+R�W!"���!�6�5sĿS<Y�3��P�]����w��`�0r��
��DF^?�����(jᤂ�dw�yH�Ja�A�O],ӄmJ�,����0��]��.�=�iH��M N�ϞZ��f�����r'eS2�e�9�	:_�e{��R5סCm|�~�Xs���(�C�I�x)�d�3Ns;�Ȱ��FAc��_��bm)��w�w]��z��9���g���Ja�y?ϣ#Ѱ\,��~᷂�d���*u�M�l&'<��bXu�
~hk8E���;��[�}�1�Ot�_����Q�[Bɯ$�B����`?s��h�	:IS</ۂ;��Ç�ك��t��@�5N�8!aa��!%����	���$���6��A�<Wf��8Q�[���-�Ik(��B�?��9��t�P����w�RE��P�,�ʮ�g�k�sY��V��!���Agh\��܋�QV��TZ��#��
��&�,6#��;�+�:��AG�ĖD0�]m���ޘ"�~i\u�J���hrm:m�6l���-��~܎�[Z�C���Zr.Xs��C?��:�m�v���\�p{b;�Y�Z�Y"�������:�>��KS�$�H@Nx�?��oL=�rcn�ȿv�v�8�-��f;H�%O�q�~ѓ��\�ŒQ��@-<��o��ou��J�KCB������!*¥�tzϲ-||�}�����+��E��|���/G/�����5E�Bx�f	6.��K�5��1�L��eRq���H�8��Ԡ)b+)�)H�g �@�!��I�yF*&���i�J�8�gTq$h���;c�u
xR�0�,���H{~Aw�;�Q�
B���֑����P�{i��5�N����6�.��'"?��/��~p����k����Ş����u�ξ�w<���۴%F���!������Ǻ@q�{o>h���{�j׭�����S�8����v�#!)���I����F��w����"J��+��:� ��D8�f��Co�Tq�=w��u�z�>���G�p�d�+��6�7����x�8:fa8~֯[k���7o���K�F�8V�z1�R �հ �� /��W�7>�r���� @`��$aJcL��]s��@1ȋԽkm��VµsΚ�fPU+8���2��-Rz�W(u7��`����FcG�A^;���.An�nƌZL���%Ė�����3]b+��&��|� �fL�l��́�3?s�����/^�,cQ�p
��{��Fڀ$��(\��U ���F7<+'�b������3`>Ur�4({��}��r�o�]NPx?������-��|�=���yO�V.U\3��)e�UlR��m!J���ƥ6Jҭ���3
sj��?��n}d�|~�W�ӳ UR�Qğ�E���i�mvg�����u�L�>:T.����mf�������W�ǟ��Uts	�|;�XȾl���0[A���^v�Ka���?�G����	�kQ�B�휟�)�oF�8j���~�E@U��<M d+�X�y�>ג�� H�l�~�n\�@4��~�Xx_���ᣨr����v�H�}���E�\�A�07u�٣�"0�b&�#�0>4��۶�w���a"S%������{đ��q�wv�k����`��,�0����������x�5�$E��������geQ�%�#��<ii���)��3`vc�+̃&�/5?�J� ��!M��������@a�	w�v�=D���`�����e�4�ǿ!H�!�[���"R�1�A�|�(v�2�p��}�=7*j/�-�	-���H��@���y�!���:���hI�'�e}��7��6�=�-���z�LO�ځ'{�#y��y��a	
��=��0��[�U��<B>4b+���B���x�A�ǎ�5Q�9g���89;r8�yb|�7.�g�{�My,���@_���F2Z���	۾�b����c��[��={
svȃ6{[��<i#|�U�� _�ڇ�Py�]��gن��mnv��ز�n?x�8=0���䙢��u�]yՋ|s�H,"��� j x0đM�	�x��?di1x�Æ������TPM�?}4�&�B=H9��7!D#��0�:!�kæ�c%�l�����@�k�l��aO$��Ę\-��9�Jf��a`���^Z�$ߴ@����:�%��7}�N ���b�� d;�w�G���CCX$� -�F^Z���y䅣��`�ߺ¯��n	����A+��F)�~C(0C@�
�/�q��ay.̅��YCT�O����uF��؉2YMa�J��ܰU��)b�zr-�C���E����>go�h<�a��/�@�U�����!�̟� ���P�<�g�NU�V׎]�b1��|5��#AZ�gsӁ ����
w�Q�+K��o�F�2B�Π;��+�)�N	A(c��p�Q�,F�<���)[�R�P_������oۺ+KwrȎNO�����OJ��9��߲y����/��Ns�$���vXj9��v��܀���5��l�����e��l��.xz؈�@?�X �U���۶�U�}�o�ѱxp�q�-`�&iR
�#i��?b�㏹��(V`p������!�'�?�CA�ǵ4l�|ۍH�Vؼ�J �@���ߍ, ��-w_��yA���ɼra�b����Z�x��H�lP�~`.儗�(�g��"� ����9$�)I�)���T��I�o�&8���AH���3���'��a�;�d�L��W-����@Z�����u�J&�� �E����7@��?��%Mr��~��k��� ��?����!���3�:0��"Θ ^0�MK�씌�uG�e�L�RV3/�a�d+e@U<wU����|�}����"G�ћ�^w�u��[�Rd���0ƶvݨ5֌�qT���[��� ���5�܂s�p>��͠C�3������y�u&��'��[�/����#�$�}���+���Mm�94g��k��=j��DOd�ư��watj8��h+���w��[Bɓm'<�Ԕ7}��	/�@�<O�����>������7�����U��x�Y�����-��@ H8<O�B��<3��g+��"�Lĵl$
�R:�Z���5ힻo�COl��Բf#fW���G����׾�]�<Z�T�20����Ԅq*~�"z�c	BB2�o�)/D7�Ad��H��F�5N��HT�$E��Y*j!��4Kg
�(��pPyh`���� /��#El*�k��͡
d�J����GՉ����>���9hE������"B$d� ��{�k ����_��B����a�XO�-��3�
�u0vy.)/3~��++�F�f��"L�70���Zs��G� 2����'�����=�;��,���y�� �ӷ˯x��>���֊R�ds�A����6;�̈V�W�U+�%y#{��d�>�����^��Z�����l;���W<�r+W
����gO��2���{l��=���;β��0�s66�ƾ��o���E���&�_��I[�:���Zu�֎G�M^�z�i_��F��Q鐺0����x��Ojz)l�@H<�Z�y���`S(=C��G��`q_n�]�u�ɥdU��k������ᾩ���Q�)�V5F4�[��3|�˓��≯�����UP�M�S�����T�����Vau�9)���)���q�D"T�C��	���i?��-��`R���ai��Ռ?����>�p�yS9l���i���^�g�p{�rL��F�V��)g�4D�[j[`�� %K+Ax���)�.Ps���N�����ξD�C���Ʌ�w ��H(������.���<��"s��!ӟ�Tu-���H�vl9h	��%Z�iI�?��ʖpO�3Ʒ��Q�Wݏ>��(�@8K�h�/�>�-�~#��I��<�e��W����0���w��{~���s��;�|�^b� �0g��@|��p>�v�eW��݀A��@?#���/}���_ז�P�����-�S�ֺ�폎�I���l^6�E]l�u��9;K Ҽcmn$�t\��$k>C��lⷿ����t����jc�[���o ���d�%��qVZ$�`�c65��L!+��-0���{0x��y2�h��-���k�Xz���p�qGc3C�f����Z��	���F�����!L���<@`�/�\�t_�B(���hi}U1gɨ�ajt_v�d>�V�z��`��Щ�������ijo�zB ���M�M\X3c��)����x��|x���<����%h�w �5�ɳ?��O!`���{�����+�3�:ׁ�C�!�h�q��ٻhPt��|�рphh�|�f���rb��>���_�^D�	��D�zZ�|����<p�9d��4�ݤ~���.�S�}C�!!��J���0��/p)��$���������|��a����_���-�ܵ��5�����2`Y�J|p�}#st )h5c�1���������h��:����7?_��x�v?��}�߿�v|d43�M��$��O]���N�����	���#	pPq9�GZ��_x���� y�J�ݖ���_�5,"y����A�}r�3�T6���_�MsU��[�!�܀- 	��i$�N��,��=�q8D^:H�H�ܧ���ڇ/djoJ,i�Xq��P�t�P5�����9������,����RJ����
�������b���]���d��F�	?��s�q/*���9���n�!���ј�Ӂ�	��0�o}�[�>��@�T���@$��e�<���<�Ϙ3�@��<%~|��0����m�>���o���<�,T�JB �g��Ә+�=�va\.�7��wF�^��=" բ<�A=H���Ʒ�F��uߧ}�Z��@P�]F�1v��_�_��~����(@�g�g�D}RT��cM����;�~Ͼ��[��`�w�3�y�B�A�~؞x��� ��'��rWЅ���C�?����QJb�:����&�`�>�s���\�&G�T�M��o��$d�H��ˠ�$��H�HLHe
�`��y(+d7�K�0�з�vچM6;w8�;���Tp[>���+�,y�k���^��(�'_~�����W�jw��N'���d�|���$?�Y�zQ��?�;�`��.UJJ�f���V�y?X5�1��H�iV��I+��@0ހ�0��� �!�z�_�NEf��yF��i Ҵ�r&�њ~\���\p7�̃�} n�� 8,NhG��U^�����}�<,���F̃
��{���T��Y�����_Q�i-
e>�[���
�×�I��{�5i�*��r�`�%A^*���%L]X�ny��9��zιچ����ѽ�������-�:.,�m�M�؍??�`�\���GJ�C�Ё!���M8�gl$�RΆ��8 ��R��F.�^�crk�0�'���}Z��s�V�\I��v⛷�!*`�<�l�NW"���A�'��z���| ³�9{�k_c?��{�U�q5�|!��L��Ar�4��ԋc8vQB�{�"�JC�q۸aKP'��X<&9���k�{)Q��د F�=�2��G�w�t8�O��?��/��s����{�<���v?�ֽ�E��?j\~�3��P�E?�B�^�Cب$0Ta0i���A��N{�e9)4�t�s��t�0�2�ʯ?��&��'���^{�΄xv���(+k~���p~������u׸0	��+Ulnf֦'��?�
������;��soz�y���/{�;��5���R�.����4׿`(E��9�ŰR��bR~����Zנ9CH#������,;m'�B�K]S)Y��|�����sA�:g��߸�=|:n(�sO퉖��6 GyF�0Tj�Ԣ(�Ja���c�q���ȜH{!y�sWo��`��sG:Y_�8��u�s�棞\�n#h�=+)�<�*|'<��*��R�ۖ�< ��7�������"�}�tM"@��#��
��:��Kv�X���Ar��q������"щͥ�h@jogѦ�7M!�R� B���1�~�����ʴ	�La�O����Z�]Z�\�
&�'D���P����*�U�&L����	J�z ��|8���Z�x"��5�,�f@���ۉ�	GNSU�,$z�w\f��q�N���;I�����g�����M� ~r7A>9;�{����TԆ�����B�Q��%,��[��'h��k���b��ҡ�\�RB�+t�#M�j�
ԔP�����۹��.�b��9U�}�������mQZY�EF4{���#������w��!�w`�$UEH䝣w,�:64��
�p���t�q������L���=�W�L�`؃>C� ���z`��4ߗ�+0�Ft,FDy�H2^v~���]�ΡZ+7��g�k"�\�;6����3��#��3������F��)"��n<�u�!aT��S6��
b�Y�<0"�C%gx9D^�00
�h>��3�A��Nޖ�ow��T�b�� �i5�iz"����l|�tX�u�+�=yȓK�&��z�U�.$)�Cl��[,��ڮ~�����+p>	i��5���c��=��l/q��V�'�	_`I�;�x�V��p���\}�cӶb�u��!�$�S��S��I��x$�
�Z���_�B����=�Vn2|��+����O��r0s�T��SЄl$�z��?(& R�ŝ�.>�&����&���G}�:�$L|�B�f������O��HS+MAƋ�ϻa x~!$ +��\|��/�4}�7Z� o��峂E<15C4 �ߵ���m���)%J��R1�0̑�#Vܷ�6���6b#k�ݘ�̗��A������Gr�T!�ԾM�4��*���qg���V|�O���\�rZ�4�*�*q������+xBը�3/�(�5MӪ�J�<�n�������=V��
.�P6[��s80(��
̢m�����ʃ��̻K'�+�B$�~M����J�P�Ӡ���ru��M��V�&�=-+)�1~�S�{h�N*wG(�N~i�"����Q�$d��]i!t���1�g�����!�4 ŀ�]� Oa��y���7�_���o�t���N�Ȗĉ���j��ٓ�r�������u�6�E^�q�}�8B[����p�����mG�J��jZ�+x�����m��I�5�-��޶ԋD��K���t>$]��<$$��`���\"�z�H�0Vmn��~�d'�y9:L�8E�0$r��<_I��X��c-��@�d������=���2p��VjE4��DL!�Z.�YZ��\W���ؽG�f����!u�@�U�K_W���Y�HN���i�g0FEz��k��%�IWM>LHbh��0ϐ�41e,=բg4�Z���px�N���x5k��o�38bs�i/��C	E?�H���`m�s�s�+Pp�m�A���~�	R[M;�u\M<q%�+�E�_���(:+O�]>�*�-���I�4a������?���\ j�	+H�5��0��b;��t�d/��uJ��!��k�@��-��iv	P��ޗ������.3M��p�r$"t҆�Ҽ8+51NͯR�^pt�,��ȴ&����LS�5a��GYYaH$$�xs��"%����"�a�J��E_�R�UeA��Q%2�gb'o�jQݞ���A�G$.,���P{?�z0<�H�{)����T�+0����ƂI "Ÿ�|��Śq}�d���=j�� �!w�=�1��l�_����?7�����vq�*cq8#l�\ڌT�M��$�*Ǐ2=�Z�4F`%�*� -ō�v�el�dÕ��$���F���6�U83ӳAI
?��Ē��V�9%]��%b�������@ɾ!C�r�H�#�m#WB�C��[IЋ<md3P�v�B�Xk&�Hާ<@b ����$�9�v�
`�$e��+6D����������j��N�&AFn��ߒh�Å?<b��~g �5'ؕ�׿.�x����]�/_tXO��D��|�U�����,Ы�A{���D����K���^e��TX�=y��'�9�_�è2*|;����(����cc1hfzzƯ��"
u4���`Iz��O	�
�N�`~f��w/���$��m�}��wY�Q'l�V݉?Iܦ��V��(�V��%��2�����?{|V����� �:�҂䛾��%>�)��Y�J�����vi��
^i��C��u_��O����`���=���Dwzf�/xL�.5"�܄uMZ'���=�Y�s�r%�ڹX�qdl�|U�ȉU4��n��,PP,�S���i6cpY������������Ҧݽ��w$/��^ӑD���y�7�Ʃ@�d�	O�;�)�^��C<U���g�s�:�FFǭ�P�#A�{�὞��۾��݅k��H��+zR��P4)yO�Y�������U¦��29{#��byh�3��N7챃�V]h�T�(��V�+���]iW�טSb�B9��k��Ȩz��jO��ǟ}��J7�,I<�j 6��Mw�P���oqfn��5�]��O��aÒg�`��H�7�C&c�����Od�cCn�y�[~���B�]8�k\�)��'�
���ύ����$���B��֬�Ds3s���cl20����ƀ=i���N�d-�2�	?�Ǘ�>
?;�>�xW��S�n�/��]~�v��A���K�/���4��
]����`�dt�_\�E���na�Hl�tNۢ��i[�U\�y�G�N���U����;<56���1�!5�۱�Ѡ����)��j+����S�O�w��%ҔN-O�'���Y�EϋB���Yg���m۶%�Ջ���!��9'�F'0�3�\:<kÕ	�K��+�3�,�w�K�/�}�C��L�#��!�I���{�� ��fi��3�lu�����);K��k�(4;�o���Z����j����)[����� �/��\��>�����]#l�:���h�T)Lz�"��ٺ��ڦ�6xpɸ���|%���7�t�둵��E��"�*�n�N3t���C�BP]�^l&o��ݲѱ���uWu�T�fe��"�?}ih��(<<M� ����+��jA[��O��o�|��%�L�����\��᜔����yخC�q�����G&�����\��0⮝Ĳ���l
�D��Q i�3M]�r�'�}�G�񩐓\}_��W�}dk-�"�E�!��l�zz`L[����rm$©O~�N|�?��@6D{��?a�#�dW��S;�������q�0p�g=�6>����Nد���{��'WA��{��^_�`7�s�N��_�e�5'E .}^�7�@HS���FU-@�Hi6h%*�%����s �'�-�������0���I�"���*F���T�[s����ک֧-c ���O�<V�˓�$\�-x����CONNۚ��6::�I�<-J�-����b��b������zh��>�������)�&�lg��L��5��}s8�s6��}{w{j��{���wv����3�+v�gۛ��3�����T��z����G+���2�F)}̉�m�= �nn�ff��;��O��������;�ܽ�v�=v��/�ˮx�5k��!���h�#�l�$�"������?��/�c`�t#K����]��g���v;p`�x|�MO�Y��iFEIڎ���A��p|i 2<���(�S�	JS��%���}��j����	�G�,d���o�6q��������z�*��@X�٥�=�ʕ1��j�A���Hު�Bb�����E�%����vw��l7�3?�3.����ܛ���%/y��:�L��$�i�����曾���,�p�n��[�v�z���v�}�:u���կy�}�3�q&4T����}�|;yO\���K.��Nߴ)l8q��s�MO��O�6O�7��2f����_��?8m��ɟv�<�iH�7�LyB��_�Wx`�?��?9�ă�҂TA��y�ۋPJ��߅Џ����n#;Ƭ�+[c�aL/<ݦ�o��Ҍg>̼Iq�����2�k-����ׯ_�M�G�ŵQ�g���?ӌ���_m5�S�T[�en�� ���'���ݠ�E[0'�F1�jں��v�E�:�Ǹ[,��-[�Q�
-e�(s]�`�5C,I	��N������&ug?F�׺g��/�T<+מ�C�=���vn����v�Y>�n�_��z�|�]��gYex��=w��w�9��[o?��;�ߖ�eY�� �w�9�������~sP�6�y�������q��yN�`�n���l���<����Co��%������~��=Ϸj��+H8���˗���rVϼ���#�i�U�]��:Y�x��+x7X��Wng���Ă��O���al�K��O����P����D�"����$#li�k=�T;Վ��׿��;��<���h�b.���7�5�ގiN��6��;�!Y��?����:��I����|�����{��p/��~�4�=��kҝ�|�@�����پ}{=�y�w���G\��ʗ�����}Ǩ?w׎3��;�<��;��?�C}� �E�۹ABŐK��G�c�6���[�G�]Dܻ���1�H��qr�?��+|s\p����o��B�F*öo�#�W��'�#��^|O���U2���}���X�QQgG�qQ����;X��X���y<��@L~�B���/��W���7n<� x#�g���t��RGS��ޜ�P�R��Ơ�S�Q�������)���U�:Ћ�NS���R�S��K�'_Fp�U�ߧe(�q=�+`KcS�ԗt܊9�8U4F��\i_���VAy	i���K���{�0�]1��$�-E�g�]o�]_���!M�R<���)�{����x�����FYG�N8�`���-Y��F��~���'7jYs��~ʮ��s����w<�~�g��fP����
��D֭Y�$�y��]�ن��lٲ&m�6_������7�j�-�����i���V�Pz�}c�\�R�tϯ���Ŀo�K0~��o��a��}��y��m[��������n;q!��������o��o��s�d���q�ڵ���N?ɿ��� -Tgڡ#���U2�p�dxdµ�4�9�L�D�Q�����PM�1���o�#��}���چ��tɪeL�)��C_S�_DB�S��X��mpe=��V��-ՙ[��{�oH@EXD��h]I�����ا�`s�*�w
��whR���+�9H�$���`9�+�\I�y�{�1��d��4��]j��zi�)Q!s Ƣ@4�W���[�S�I�и�GR�b�$��3�-%|-�豸�Z�1�l7ݦ�Y۰q��E���	`�;G��ƈ���6]�-����� �R���zd}���&����w�<��mXw�{��fBok.���M/�[ȕ�H�=w�m?��W{��*�Ɲ�w�b�y��v��N�d����XU�K�e�����AL�Ng)��г}�ͫ��!��0���P�|����M7�@�\��?�zB�c[t�l���=67�f��#G��<'���I7�E͉<�}�o�o~����ZǦ��m�HSɑ�BL(F�}�V{�������	�KlzpP��L*��L�k��"h�LQV��T�Y�.�g�E]��p�&���̝b,��k*ً���J��q�͈HZL��k|�Li&iD/M�O�h����x��� A�&02��5��B�T�Q��<VR/�TkH�N��1����7Xn� j@����h��5_Ms���'gё�Dl��}b�<R>SWg��᣶���m<:��5�Ǖ�
�7�%Y��esl,F��x�nإl#�?s����^�B�LL^9�8<S	���Ӏ�����`Lh8DB� p"dAspG'�"Li�R�r�'��e�(lT�c�ר7|qt�I��l��hZ,��TԴ�js�Te���{���[n����]WP���fQ�vO��g-��ZN����:��)T����(�ry��<L̉���� /$�|��y����H��d."N_qW}����Z�n��!���<� $�RB��M	�E8���ko*���I��N��4'��X�����ԝ&RK�r�W�%MC�!e
),���1�=�\��z�l�E�b�������� $'f��	��>����^�֐��]bip��A�RoTAEiiG�=e�;�:M�N~Xiv�V�]5�o���/�|�ݓR�M�W���B��ֽP{܏e���ZexT��4/���+?��#�#�c��9J���p~p�云�1��83�%�R#�Sw�6O1!M
B�u��9.��lxP��'��i�R�#�:b��G\Z����uu1HC�l�m$�[��Vk̅��݃�f�N�L ��}�s~ )��я~ԋt �����A��v�o*6�b��Z�0�9�	kRM)l�E�6O`R��3����,�v����Z���~�C�f!ց������)/�ą��`�}I׸Ѧi-B"����酂t����m��B4Io�1����N�s%�J*�4-b&��S%u����MꛘIJt�0oiM��_f�#�Ҷ`+����]�D�G�$~ER;�'�j 
*�I���<(��>�K学��Ms &�{5#����2�*�Ij[-��\��z\n�|��*�z�o3�?Vm���p���̡D���I�@/�������Jս�0���g��?�^���\;�0w����m:}K���@V����"i�7n8�?ɮ���c���K�4�{�C�	O����(�b�*�/�����a��g���a7���xҬ	� 'ok�֨�C�<b��[�T�3t�Dx��Xt<f��Q��~ac���\:TIWS��h��S��d±�y�c�
�]��6��Q�cY�T�f3��ii���`��}�K_r/ ��W��U����&�w�Pe����J�]�����T�?H��6R���C��ߒ��{H�ZYkŜ+�j�7ˈ*$�H嚛�r3����G�eҤz%��1N�2'1�h���~�.�`���UW]խ��/����uBJ�L�((�)�EED^k'����:i.S��bAz�$5�ߩ�Ͽy�~`��I���٠��-�l�t+�Dx��O�.E���ͯyJgR?��x�N;��	;p�q_?�w�w�%�������1�o}�[. ���o�׽�u��4^i���K/��|��#���5�"��g�T�u�6;�z�ӂ���iB�/��밖-ըV�Nx�?����k�,xp��]jc#�b�G��l�c�mzf���IĂ���Gm���v����!����&�j��w��~�w~� �R6��H[06� ))�F�֢�I�g�B;��KʡO������!��Q�����a�b�v���p����GV�č����
cÞ��s�׀�$127�Œ��\�P��Qaih|ǵ�G��Ԉ��#|]7���o�%�{!xz��J����E?d���r�|=�S�O�+���`v��u��������������g0~��7��>I���h(���d/�� �J|Ιgx�D���%H�h�A�i�,A]���>BK
ӉQ��@�觠4�*R�+���;�Rږ<���է�^�Do��p:��"G���O[����'�l8��k��f3��2�g��U�f\Pr�𑊯K�:���^W�o9�1����Z�?4 #����m����{�Vu�"��g:���6w���5�,�5���k��Bb'>��dtc"!ި��}�s,$��7o��[ny"0���P��DKk���?�.}Ƴl۶���1(P�߯l lr�5�4��<h���җ��Ŕ��2$��C��������=?d�F�8�p�5'���Ӟt�8�� �>�|�x"�M0n�'��D�&����F�ĀM�
��� �,�k9�h<HFƆ&�!๤��`2_�.���H��@8a��%!�-�l��!A���]|�Ů�+�"̞���w뭷v��@�!>0<�R�qE�h�It4�����A�!�`�3sG?��O/��wa8�^�>�����b#���@���x�'�42?ϔ��{��W�H柹�H�x L|Ƽ���\�#&s��A�b��ꓰ�ZJS�N�0w��&I?�S��A�EO��Ko�f���!.j�x��pK-��?g�N�jW\~i83hay�T�ߛ�eU2�ļ����3c2pb4�����e��A�0Rh�'���a��O��w��q�96_mط��M;x�q����Ex��v�%�k��,n�Z�;�;��^O�r<e^Nx�?����G������U��~����g_ye��Sv��ٶg�#{�ə�y��~#\x���áYX�S����1|��_����.���ȒhW6��5�yM�����Յ�-�����;ǼH�R!˴i��G�.�wo���^0�Xp:Q*,"� !�^�
c��"������5�saTC�s��0��I�A��������"9qX�~�p��< ��%X66`'y� ������Յhn�
qހ���?��3gR��ŕ��<�	.��ox�"am �H��ƚ2<��t\��[�������#���1?�@<��y6��y�X��w�ß�e�!в� �0�J+��z����H?���v���B�w�O�k�����ؙDj��Q�`r����=��nl0"����#�´��5�����9F�Zj�Z�	`�3`���;��EO;;G՘��J�8{��N��w�+~�5��.��מ�c&����?��.�ǚ�ߘOՕ�f�\��0`���c����]g�sٱ.���m:�p�+�a��kk�m�����H�n��˩
:��ۊg�N򖺖�0H]_���H
�2T�3w�gO��{�F٨�����t�MN(�"/!#��g>��@��90��]����)L��r�pl�E�ߴ�Pζ����*�@���ߎ�����+�(>$���VaqK��vߧ���o��*t�&O���
�8C��$^��A��;�⁔L�(BdyLAFK�ć�a <��z�R��?���l���BX����ε<��5��v��F��Y#�0DBȻ �Kpu8D���BZG��`\ya<���0��������\3��O�`2�����D��HPP�l*�Ë��H��^�җz?���Aq�����{�0�fO��y.�/���ó���jg^�/�m�� `�E����Fgh��"L��+���6�����Y�����A󥆯kP�6�`tl��ȯ7�\�/ʈ�%{��Tm�V�9?�N8t��Y�.�I^Br��������������~�;cK�N��g�3�v��}��b�]�%g���Z����O���1�+�aܴ�Ȑ=��>����j߻�6{ы^�O��G��9�g�a��c7�tC8��,I� ���w��UY�j��s?�sV��!�*�� ��QX�b�= A}��a�MR�uLK�(����V���A��s��˭��ѱ�OYA�ѹ�)o��֬�����F�5}R>s!� �8Iud����XUm�[Pb�D	�n��B�!��`y�C�3!�H�D'C����P"�qߣ���2�;#�N����!�2�)]8G:r���C��L߸��>�9�&3�0J�DzN��p�Xb���s��	�M�%�^�s�0�7�=�C������ɷ_�s�b�g<���	k�>��^<�x/ϓ��o�2��I�	�b�0��K��cXZA������vػ���;h�A�m Q�2b?���zw��w�c4�GZʾܰ!B{�G�7�}��Ky96�x��}�S��=�G^`�}�U~��:� ��e�Ұ�����/	�Ď19=h�Hē��q��A_��t0٬D����|SOL�q)��٨���Y��h2�	��|��ԧ>�Ź9���/����!X�WR�F[�7�����4f\M�b��P�e��@�[C/�\?Nl�O��6���B�|持��Ƈ�-�1C�������i�E�Q��q�H� �����ġ��sИ7��?�Y;�c�c.!�<�����!yq8a
4�H?�Fy'k!�O~+�C���x��$�2E`ƉF�{H�"��i�f �<�>\{��A���5h��E�1a'A��11�J���0*ր~ ��,	$"<�*#3sGc��H���a ����z a�AE0C��z�C�!�\#{�y&��z3_�����1�^�g���y�1��D�4��=���RD�S����΃�8;�By��]=��X7[� Ͻg?�*_'�L��g�9��=	�O�T���xff�v����n����Ӄ���Y��F�<��Y\�"��flx��t9�?��~߳�D󲯔��=;�+�y���^��9{$��#�_t�i%s�Ң
ד�&F9n���F�!��� �>�tH叾옺x}�vl??�3�67e<t�>�ߋ��ƭ�A>k�"����i-Vي��ϟ ,I���!��������!�G��F�c�:$Y5{��$�#�qCp�	`�=ćk!�ZS�!}�A�a�H��%D�y���_����� �a]Xs�v �:�4�OZ	?@9����!&̌�A�!�"���7Z��A�Ȣ%HC�9���� 0�����|���<m�Ly70�"M�^��k!��+���yd 8�Q%�A��}%+c��,����� ��|�o��~c,�V�j$�Ѱ�ܧ=���4�����4z/ۘe��y���u�].���gنM۬2<�I�b/#�gj��+:=2�| ��q��o��k{�A�!�1��)F�zMI��~�)�`����>�/0�=Q;�d���5������(�,Wm~n�\�s''��t�B��j1���/���
G��� wN��������Un_<��a�(�9_@9����u��D���kn��X��H2T��Ѣ�]�ɦ�v�7﹉���7<,�#�Qp���6z��J�Æ�@@88�D��o���Ɗ��R~��4\;-�.�7wfȔ߹����bǏ�R}����ɯ^��I��=H�rߤ��4�X;�ʡ�����s���> �L��&O��B�e`�/�[�ϣ�a�`��H��	s���p�>6�'����8`H�M��ɘ��O���y�x7��0�`5/�$�����\9�3Ew+e����@�����r>�qu��b���bzs~
���s�-�	����
�w=_�s�G;����ԟ
C��>���0/֗�����U��4'y��Cl�!ڂvkC�[���ͷ;�w;��ʼ�|v;���saP!X$r�,�c�Ĺ��&o�}���R	�$|�vb�W�h�4F�_��_�_��_w�3�� )�.�_wBɁH7��4���6:��B��!�p<���hƒ/e�7�"�|���4�q�����%��0u$�P!6V$b�{�l<gy���&�<宙F��^�S������C� ~��ȍPy��8$qy��7����lt��o���~����l<1�5�
L#�%	�@*��TiO��f>%,C"?�ٲ�X#��wA�h�B#A����G3�Y�xJK�z�4!}��ZZ�����$Qk�5W\�����8�vC[��J{��-�xK���.��ՊkQ.���z�������u2�	�ŹG�VW���cǝ�9C b_)c�������,h%��w�P���S'��-���\�K�nl��|;$�%�˝r����+��.^��|�qCG8�������A--�Ghg��)
Q��7�#p�x�B��</���p�W�Y�%Q��W��8D��`�N&DCɺn��B$0�}�E��d3(7��i~������o�I{�{�c��G����R�$u�ͽ��T���b�NAW���{�*`2��s�/��*	Sp^%�:�|�HV%HS����yz�,W;��
�V`��1�*xP�RF������� $��Rp}�s���� �Zl`�@�D��adozӛ���4��3�O����f��I{�A^\#�V�z¨�c:�2�k��'��	��0V���}���|ݫv5�5'�@����S��BA9�b�.@i�n3Ȝ�3cD�~P�.�!Q�����A]��ix
�ت7�}���2�6�n�DD*�?��So;	��V*��({����B�|'���R�ͥ�\њ5��� ����z�U8$�T�����ẇ�k���~w��˳GH���E6�.�K"�px�T�:b��W��'�nY�`�R�s���L۝�H�TAD��0p{��{�ԩ�5�D�%M��Hʥɏ;M�JҊh)���4�l*zF��&��RI�&��&`CW��O>��VD����oi�`�A��-f��c�g�)��h��]ஊt�D����ް��w�>1=��T�M��2"��U��[�-%���_o�~n��-�)�c[��3�/0�@�9����p����~��ֶ�y��M�f{�c6ng�n3˻&�7�F3��U���� cFg1O�W��񮶃���张̢0E��R��e��CY!�N���2�b!~��V��ϧ�+�\�&��Ri�Z�Z�v.&�r�' ���B&M�,Ҍ�:"N�p�5��:�{�����?l䃇��Ƀ67{ت�S���RD�$��v��5,�)d�I[K���?�%�J��Y`�TAT����q���H�H����C��xC�O�囘� �x�=���E�щܐ�	���&?�7ݣ흤�D��/4lt|��v��*hxl�S:S�	�A��k�-�BSFtN��i�i���\�f@�C����w��#��Q𿛭�f�t�
O�v�$5�jC�Q"m�W��w`�O�V��b��XʱPT*��E�)%y��3('�6-5�*�w9�Qj�l��8���x��c�Xo�@�|� �/dϴ���$��9��)#'������ϵ��q�?��=1�����sI������~���o��0��1�H�T���[;&v˵�-aM�%f�g�=�����5/�a�Uv�}�&�gl�m�7F���kڙF�g�`K5i3�UE���������vF��Eo�J	���\����^�|�[�J���d� $��m��A����S�q@�C�OE�e����� -2��S�JM�y��;���}���{S�}+��V��sso��9�����k���n�bwio�ji�I߽�_�w{��٢!(�8� ���=�y�8�Ѳiy6A�u~�l1���g������ ���o�׎?ꖂ@�y��`o��2"�ԭ�x.\y�%>c�����,b�CS�y���t(�"xMj!�C���� ��$E��ԷS���(9�QMk4�b��?�JX(��F�.��U�U�<���^z1w�d7�HǆJq�w2H�c%k4���)�.#F���2{_5�q�8/�Kl��٠�F�c.�[�,�1�[��[¿���{r��{��l��7��1�胱��-���/|ZU�jH(*-3m�F��m.mBY|��ִ�����1���w���ش���5t2W�mgƎ>�@�1����x9W��C���p�F(���K=�۟�7��(J���=J�
�5��}�m����(�!C���H��t�8��B�^o��C�l�S'-�rm��6��=�l߁63�g:�X��ke���BZMk���a�-�6�e�f .5�[/W0���؍��>�Ϊ�1KY\����l��_w��h�:��V ��*^� �8b���.*}�LF
��C0��'UX�s�=ç9㔰P:C�i6\�ѩ�C���J���{�z7kh��K�t�ދGB��&�W �e#^�R)2��Gy�i@��c����<��o?RlyY)=�S)������x��V��xtσ֜���Y��#�{�68�4
��c�`��h��9�i4�jQ�ˣO��c���֑bX� L�3zx�B.�(���p]O��f�GP�L���)�8��ӛ���pH�Y J�І���u��q�6z����\8��H���=���<?o�*�k���$ɷF�:ַ��M�ۻ�����gN�sAX�mf�4�jA1�4(1}l��u��l���^<i�A�GDe��l�m��Yrɹ��+��t�b���S��!�I+!AB_�~���X�ݳx84ۊEu#�a�U�ޖ��.x4b��ʵv�78�?¿X�� \�ctXO]�fpl�Zq����e@�H?�W�ݣC�v����ڵ��l	�DؿȔ}���:~���QF��l)�xQf�g���w�7;�9�(���[��thb����@��P/FF�o�s���դ)r��W�RC�9�R`J�y�K�q���_�u�Ycf2X'eg�t�C�+�q߾�v��;���	+v+1w8�~�3T0Js�(FEX�mW�
������� T{0;?��� d�H��9)��;;��-�'Y�m��Mv�5��=��a�y�aC�5�޼�;�o�s]O�hw��ʷ��O��Wz-P�����W��I��~R�N�_��_w&�^�9�?ˮ��*۲ꐚW ǽ�p���;wy<�{��.���ډ3�+v���x<��z�>e��,�x���꫟f/�����#�7�b��N?A�5:u�t�F��M�(`-$ �!%�L 	w^G�� �����5���^¿ ^9i���A.�?iǚs*!�m,�ȩ��SA���S�D ���}���g
R������?�`8C�sJ�¡��-���6�*�v-�5�d�<=���`��V�����1���E?�9�I�����2kU8_��ʏ����W��X%��9n�	�Xj��߲ҕ���	�ѽWE�O1(UO�ޫHOך>�����T��Y=c���2�^�:lB/�b9X�e
9�� h�M�c�a�XS�x�b"����V���&$=��/���e=c����y���ʯ��i�c��q{�w�]�4z.�����0�i/Ɯ����aՒ]v�v�,�`�o�����OkI�EO�%�Y/��/K��i5���`�o��K^�"p"�v{����o���M���~����.��R[�f�5�mgy�RH�*Q� �P<7}�o�[�3h���^+�����"^�q�	�L}&,Jf�y��۴����=웶������8
����t���Z6"H�� ��Vo�TA�f�k�8m�"�Q	c�$�T���u�W�Jx��ƙ/sRe�)ǉy�Ŝo�!���L\Li1��sD�s�񚠕4Q@<>\�^^�x~�)#Jկ���� .C�E��1�7�4����ž��(w��n�����7��Iqn4fmr�v�jC��-Y
mv;�,ve�k�f�s�&����f�n�F�4�������3�8�c�%;�԰��:���S'�ѕg
/���p���k�pf ք�si"��9j�zw(w�;lF�ú5k�&��z���Лv����W�h���u;~���DXl�w�];�ˮ�:�k79.�u�۱#G�?!�b�r
7^���|�+_��n}�m�h�������Nu,���!�=��]�a������lf�D�\:��6���OeHx���={���g��>�����݅�;�����pg���V���n�
ȕ�W�]��x*P�P`��<��g>�Y'�b�_��BO5U{C�!�̙�1�&('x:<g�X�����wZaxpD�FM�g��5r\|膁渖ok����"(�����4u1?Xo�������q쑱Q_�:?���D��A��uk�z�0�����gW@w���p�T�)�߅bֱ������ׂY�z�:[�bC�#I���Q	�:��kϟCDn��0��a�Řbm.J+�e�8��m���{���ҿ��;��!U�q�5��u7��T3�^z�S~�C��1�J)M 9��_잣�O/˟��Y*XU͸�ᡟ�:IbU�����^5j�.X�<:�z���C��׾����v���C��!��WJ��>��hr�0<(�U~�'^�^	���C_�<X)�ël��~��{�}v8,".��N�F���cq�g��i� Z�<6@���kEB��B�@���?��@3 m3��=z�K^����@�c5!�9��P(T,u���a� ��)�a�y9���պPMVd53W�)�!_�� �Ie�o���qm(+<<8͕ J��v���p��;�A^m���C`p?FǆGFI��������X�Pf����7����\8�ڱm�Si0w�k��͚R��<�_o)*��d�cࣣ+m3m��(�f���n,�,,��0$`�Ϭ���W�Q$cH-�'���>�g�� 2����e�U�ׯ%<�o�sή��
��w%�F���O}�� .��i��o{5��?���v���7����/�3X�q��:��YK��_����Um�u�o�� �&�R�88¦:v�MN�� k��M.��x����8�#*`�QYs����y
Xt�z)��u����EpO���-�u� XA?p��V0���52~���;|�#��H�r���2E��X�m'����~�y�#>���ѹO|���� ����[�l��,�Ga �x&��s%���h��q�5kW9$ǳ�y�]~�����\�q|^Ûcsc��9#����(����!���k�E����-QT\J��̱yM� mjR�|)�n��5ǽC�n���Y?NW�.��Șٱj��{	�V����q7��m��I�J��P ���{�)T9P��s^�a�7rl�F
=��]�z��q�����=��ɣ��r1��k�s�3M/���b�䄑X���������.��a��+��w�;�����/���gݶekx�-k�j�#��7^ikVӏv�ff��=�`eWmo��4� �og��+M==y�~���E�B~N�K��K�sW��)q�b.�^����j�����>�KG<b1/}��Kv1�VӨ)����'%KU�(�#�Dt&FL�����-�"����/ӿ��Ω"�p���J�yFT�JC4'������;Ne2BQ�Xxfs��~L�;׆���t���N�^���nܜ�&�0�3�=2=x�(
Un�lX�^tA @����}�QkD�+�{3J�/�>;���ZA` ,/<��銻}��6;q�S�[(D"8h���aO��ۥ#v�nŘ�O])��)���;��k�u�4g�A�¡ D��*>�z���Ԥ=��=�rŰ������#���v�G�R*ة'��ذ�B��}op^���z�g� �z�_��Rtv���XN��� �N�,����a�@fV�F.�"��v=h�a���dP#���Q�?��?�M�Pb! U ���Xo��|_��d!(K�x�Ҋ�Ƭ�*0�6�њ���ɰ ໯�p�.gt+,��l�B�yh������]X� e��������X�,�f�����P�\;K� �5&x*J�󲱸'p�K�=���~,0��g~�g\� ��g��fR������[�ͥ�s��=�v��
�d�_6=�k��g�ry���kF�?���v%����'̕��@�̵���kc.bC�U3z��2a]�X�W�s�p>�g��1pϸ/jCyn�QH	tm1�?)�<�X�_u�W ��=yb�V��|��6�L��I�pK=���l,�6/eee1�Y�@|�4s����«{��{l��Ƿ:�g�E�p����S���0�B,���W�<��̉���?�y��IY���(��̔oڑQ6����A*�U,Kl�)��iz�f#�T�u
f~����R��y�b{!��c���9;tp���}oX��66^��k���E��@YZX�۷�#C����+A܁�@F��E���k\/��DM̱���5���N"�k������:΋@�;Vp6��c']�#�Ԝ��،��^����.3s^�zE313�XPףt\^G�)~�@�o�r繂���|��Ԁ럘��������Vf���G�P&x��ȍ�qn�w��^
־�1��	؇�T�8��i�FA�5.͖w�b�;~Ć�ﱡ�UaM�[��{��k�#���S�����
��������a�������7����z`Ȩ��Ӛ���ke�(z�d��"��"�@��b,qxd��Z�"W,O�"���)��>7��l�]]Z'���Ց�)~=��K�r��[��7l��%�V��p[�l\�����?�������\y>wki^���e�?l�sAIET�3g	��E�(�"��ur�[͠h,X����u�0����H�s���j�
V��/pKA�2�
e���~b#x�pB8��`��^�ʯ�?~��杺���[�¬1W�k���.�q������#�jժ�֨ovܡAM�/Ͻ�9. 9��ب7�n4��ޭϸ�ߓ"`�dg���}��ܺ���+"$�7�.Jx��5���O~}ܓ���%�l|�F�m����k,���~�w�r|��Wlz�7���;��B���r�����(��[�9d�<Pd���/�y=�Y�v����� EI\��0/�~AJ[M���<U��0�RC��& Ȱ�qTӡX�֧��i���TťF�!���� �뾐d�p�[����xk{k�T�e��1[��v\r��׃< #���S1hɕ��q�Q�����[�?��'��\د����ۯ�����ҋ/� �����)��JT�%�@���Q�t#�X��t-�W�@3�ylx$�g�T�K���R�y���j�W�!K;���vX��9�k�{�iG�����w�k��9�U5�E����ի^�P�0ؼd!�����j+&�Q!m^64�D���>;z����e�*��$T�˖�B����Y�g(�
�m{��^
 �}bO���0	N ��և4����pN��9�Q�/֋Z�?�wP��,&yBx�2�a�s��fD�'�+X��u|�s����C9��zZ���1����J�L�5悧!aԣ4���f~��c)5��B������.�E2o5@W<F���Ҋ�MxWR�D�K��X��� ,]JR���v��z���PŸ���R�.='N�f@�3�^��sL\����(���8y�{�T��'�Z�S��k�(_������B��~Ϟ=�'�'��׼�[���-o�,Ω&���W=ﱆQԫ׭��bSӳN�7^̮ەV���ȕ�e���Q8ݵ�Ϡ�Wp��b�7��W<88����_���pݵޡ�۞���C�e0n���uހ�߰2<Ԫ�;p̨�A����K��y���wz0\�\v�BXW]s�o~`m�٬� kyfz������f��m��a;9=���iD��r\� y�r!�+�y��~C}dU��o>?���`�"�����`��]�U5C�H�_�zsU>#��&���yO�T`�X��6���P�����>|�M�5�y��F癨Z�g�޳�_躽7l�M�1���|�P��96�������ؐȫ�[V����^�PR�Zi�8	"Yв��B�@SN��	�*ӊg�ȩ��e��U�:w���ɭ~>j�����c����W�Y�4΁�H�H%& v
���DY�z���H�W�4��eu7s��\�X뭬��@'�?��'&��|���.�](؀��2��=i�&gmhxܠsvt!�Y���7���}�+�؁�/��灂�"Y\��H���"�L�.9�Ë}߽��ϼ���Y�x�6����AV��]87���[��E���s��n8>�?b�T{F�Ӽ��O+6�!��bx������+e�ґ�>�屑!۾m��_����:x�<�a����CA��=�U���BV�������.�!m��K/w�W����&vh&\#�3B�F�@{�	��`8/�
�C	�0�xE;Q����3�u)F�2�\�36PP0�	e�<H��~��x<���o|�=���Z�(pu��N �{� g(�����q��|�����/��9��F�=�<o�d�[�� 歴����=���=�뮻|=)�V7K�˛J!��}Rn����LxJI�8��RPEw
󤰍��������+�,a��+���-��!�+� �=X{����_�����a��iZ,�g�'�{�}�^����~�����R%�ͺ-�o���@x���<P��Y�����u�:�sb �Y�x��o��M�k��|l�~�k����4�A�tl�m�y�%���M604hS�s����B����g��_  �f��j���ȋ�O|���[���m�~�w�yd�^۵�A����+H���˞f�_y�]|�����qc�k��h��_�W��y�L��E/z���%
�C8h#�z�ڂ�ynz�>��OZs��!-��1����5@�<������`��]R��+��źP���z�k_���?����� <�������T4 
�J�K"P�%������Cyb�*�&�0L���tL�/�D����gȖa�!Xو(���o��m����i��{,8Rq�\?��?�0X.�h2}ڲ�Q"�x���.8���T�F�=YK(���7��9���7�1���^ )��e��%lH��f@�Eֵ�q�P��iuu<y6�w�
l�C�N���dm��.VZg2���{ �y-���?6e*���ݳ��{����A91��-/_�6+mbr�ceP����;mF�����'�vvO)Q�C��d�Gq���+5`X7�x}�C�֭�b���>��]-W|Τ��_�=�����z�&��a����g��q�q��~�
ݚ o?˹F�>��Ϻ۲��`��ƛnJ�{��~��`�+׬���.�e�"��E� ���ᘈ�������rx��a��Y�A!�$��<��wx�w�=_����`��:�!�(�u>zl6���rh!�Se/n��>�-/�1/��Qn=�M��MДkG���6���Kγ 12�E�	�b3pl�G�V$���*����̅{I�%n/
��3��=�H���B/�����;��fnT�FOf��/ރ�Ұ�����`����VQYH̓�^k�B����O��	b�S��Ҩ�F��'� ������[ǂ�u,>�='�h�S���1�*W	qF��W,@�[�B0����Q�<C�-o�����[���ӟc��1[�r؊����ʞ�I�;�=�5�6���yn��K�o�} yld��R*�'�w�?\�!��M�X^ׅ����FQ�$���Xx��֯�U�/��n��[w��?u��2��o��6m���0�w���ѻ?����+�Y/��ֻ�;�T1p��`�~d��ٟ��^��Av���k�k���HŬ�:��X�ln�VA$
�)��`RV�\������tK�E��������w(
B����Y�Oz��T�f.;,�/��S�V_�e1  ��IDAT�9�N[ذ�������
��=��3�&�
��,|\�T����@�\#�8��1Ҥl�(�
!���Ȇ�ް�8BOE���Gys��e�f�R�����h�3�g��E�rI1rY�\�,e:�����~l��!�Y#|��B��s=��ǣ��Ul�$DdK(J Kp��K(+� ����
�+���4{DB\i��e����|����$#�y�K橸�2�4o�)-EvU���n�Ev��WS�y��V���gf���[��+lj���1�|h�X��O*���tO=#�򛜎�is�>g�췗������~��z�Z^EVpr�{�����^��^�5<�<X�+l�E�mnfֳ�FG��.�+~�#=�ȁJ����9w�8v{��O����N�� C@��Y��@,�w������n��6�,V�ɐi�,��Y��>v�G\`i��0��@����q���Y��=�x�;��X��%J�%1#E5(�JǙ;K���
E�}
��_��]gb�D��oȃA�2#�	sF���#\�����pl�9� �V�ŀ�&�{bGDx��;���?`"e�7/�����: ��6B�\z} JE�[�����r~�q)���
��X��^��;�c.̕�t���qߠd�C�,��3PSp���|��ZB9W�U�Pe�p-|�����P�fjy���R8U��"0�#�B� ��#��*��uy|(��� ���y���k�xf\� ��?�A���c����8Ć���}�T����U�"��{h�f�Vۋ�ʵj�������E��@V�u(F���5�������]D�X�y�S�[����g]��-��]���62dM0̠�����=�v��G?l����3�ckiI����6��ހ0�&�ed�<�QK����}&XjP ಣP�G�G�Gz8,��f'���k�"E� ��q6�d� (X<��ۿ���i^�R4�u]YMMUm��	+���κ���wߧ��r�c}���c�C�{���@8^x�_��}�V�QH�D��9�"�6 �S6,��������TF�
������
G�1�!����B �>�dc"�`׽��r.�P%�|�7�e����>��7��
�p�@ �!�U�P�?�˵s������b`�PM0W��'k=%����d�=��FW�X�y��,U/�kn��V��ز ���Ǽ喙0�geYO���{)���=��e8ʑs��Pp
��.�4뽖Ѧ��R������_p��l����ɪ����2͍���)��[#��s��ǗŶ�@��Ś�B�}S0&/��J�X�������͠+ŮD�r��q�����,�L7���k����` pe�{�.?PQ�9�5 ^Љ�]j���
��?�!�{��͌�˩�x��	�]�ͷ4,��dq��45�ZeC�`�������/����O��
,�3�����Mn�⡽�>,�^�V+�>��.w���-.��5d5���E�@pE���:x�+_��닻�)k��]@����`T������T����l~��jV̣��:J���	kW�+c�%��W��7�r�����ͼ��:O5D�U�&�e{`щ���'�'�G��֑��T�(�+����\���&����J�w�f�Q���hrr�_S�XP�j�Ny�"!�'�|��"x]�(3k���W�*2���L��u�
��B��_R؉������kG	����5����J��u�&[�vC�C���F�f��2Z�ڡ����=�p�IH�0եp�����T�Ǌ��=���S�>�;*ume�Vx
"����no̿�]�'�]�5�e��Q24�7>ZT��B:5�� �X>���M�<��M�Wit���k��`�u�b�F�����Nc�n����pz:����H�Q�
T
���B~��2L�`����� ,��?P,@-Ef�Nf�7i����g�0r�<�ShcJ��hKA;s�ֲ�����"!��+y��z������*|�^H8����dR�^�J�F���q}�#c�-%����*^W� �3�,87�e��=��o{�E2�����`�c�
�K��p������\熍�eW\�ﱽ��t���=�����u�����f)�<�/$,��"�U��i��vs>�薧}�+
�#�?I���_z�Vw�����g�#>\��Aq�U��ǟW�]�٨��+k�_?���Ŝ��=�=8������xj���6gJ�Y/����q�t�eeҼ��n{�MۚO�K����nXWX���z˒����K�Y
��z&+����)g�B��Uv`��� )�>�8�AX0X&���gr\�,P M�N,<�U���lp,HÁ8��9��8J`#ă/���p��b�*$��=T�
�HlŋUJ��x��z���,�� ��9�I<�(���x�9�+׎@d���/!�g�G���cP2 �Rذ�|�����ٟn���z3��7� W�UB!�V��WU��2uXlz�9�Ph����
v#��\|����s.����꠆ף �<�����j�9ǥ�u%��5_���+��ݏů�n�#��9�ei�Sa�<��=�z�Iߠ{h4;q��b@5镲 ��t���)���?�'�5�<P*ts�گ��BLKu�"�X��sc������_�a�g�-�j>�E̕@K$K����<�����))��=<,R9��~�^���yF�K��#�û�M-gF�5�"��W���^2��,�Y�W�&��{�U׸ %�K�
��I�;���{�\���Gq�7	���0J�+��Pmx����;��L}�
����h��LP4�B���rl�N)�B��CJ�� ��9�
����5��X�j�5�f�w������,���

�`�ū̚�j5� ����x���� +J���2�!��0�W������7����1�N!�̑�@�F�P�iL(BYJ�-o.b�B�F%��'���y�*�z�b&��B���S
�̯����ql���(ԭ�l)�<���B���VF���4+�LZh���U���`�n�/�p��m��gPP����c�I9) �,��^@�s�e�� �2x�E�����F����������p.\�au<_�=���l�ѱ�3x�:E6E�S������M�/]kl�"��d��ĺEp��!���۵k����w |�4W�늴J,o�K�t	*	8��c����y+�4B����_A��H�D��u��7��F�� w�X�j��2R�s�-�5s�(3���ÛA90v*��!�D_�y�����+~e�(@�5�I��$P|�&�7����hE�Y*�|xA�?���\��E��d��� �h�����Y����\}��2���,.%υg�ץ���'��f��ĜQ�<_M
�i��"�no/6�]=����Bs�p�C��U[�:�̍���9O���Պ�n�� �<G}L����5������T�d���h:��E���0�b�9Z���?�������9��3Y8< ϭ.ƻ�ng<&����Sˀ�|`2D�'#b3w��  �c�%�=�J�;q���}Ȏ���
V!V6OS��-�O'��S�TQ*X �4�a����Z�H�!@����4]EFlz�� .}>�1�TʒM�<��s?e2�F�qQ8X�X� U_^��\�x�;�ax��L
#�J-�\��5�=�X�y`=��B��� �a>QAY�YLɬ vz�h�z�:Jc�+u%���c�O��&��5 'I!��<A�xR�>���m�>�_1Y�xO�o�פ�Vz��I�H��!�J=���N^���w~�b�b[�Jl{X�1��	*����.�r�_#�V#��Y+-��n�'U���Ih����x@�qnJՍ��R��]�օ�g":����3�.�g���������6`NY�-��}ou������W�7��).o_�5�$ L���m��p
k����c�lr☍��j�#�2�}��+͔�gyZ�!��<�����o�'m���%s�_�`�>��Kإ�����"l��:�G>x@-�!�!�KU���e��"�
���!��+���%��2��`05������ �X����=�n]*fJy��kd�xR^�zRПav����L��!��)K���K��Q��k(t�T����������ͣ�"�w���3n�նl�(�����~�a]�ךd.ɂ-'�l)*��g��]����������9���٨ (ҀX�N��)���nVx�S;Ik�">ǉ��{[��	߲��4��h�W$ռ�Q�h�~�w�x�2:a^�v�;�6�E��_7�s�ȫ7��r2��S4[u��|�U�q����NA�,�>���i��$�ѣlwb�03�T��5����A,���p^]y�l"��XlY}���V�v��c��J){Eo!,�f�b���=��٘�e���@�|A#�a�#���������6� �p=�{ѵ�]V
!&]τ�c}�#OP% FL= ��e ����Е)�Fձh��|�ǀ@�~S? U��ൠ����|AF���I� �@m�><M���L�Ac��&hG�>ץ�]�,�@x��s��f�(0�BF��f)\���0�fI	��N��Z�����ܴ�����~�ɩS.\f��5W*�zZ\�
p]k��n��sn���W��� H=)6�Ou�4%��$:����t�3���m;?W̕+�
��O���^~���-W�P%�ً��'B
u����=/�?35�ߋf���������-��{����F*��-pE�9wP&���t�)���9�X���x}��۹<
���k9�D������4#L.ndi�ܞ�8�F�"��z-���*���)>����^B?��+=u=a=zd"X�E��� h�5�A67\�z��Y(s��7�6�(��SgScR��,0	8��.X��M������0{捀U����P�g�����d���je� ���̊���s`�@7���~���>�<��96��<,w	@��T�)m����A�)�ϛ���R�����86�'�+�WZ�80��ԪR9�R�R��$,w\�.*�ytM�:��w���o�-�̇�������yC�c)���3�"D�\�=�}��
�����kIXCs����y�
r�6@���	�[z�L��,jf6x/��%��9/جt�г٘�}�w�Z����>׾��1sϫ���(dJv�R��f����7F�e�s��'O�c���#p���-,h��N	�c��Z�:�?����oΝ��;W����nӘ��3\���2F�%�.h��\�^5k�*?l�Us>t����e' א�'�[A1Ǣ�D��t�?�͖��x��a�
�xF�\*����U6[��M����d����[x��s��s!��p�4��5��'Rl�G*]/~�	�� �W.�R�<�e�I��}��bl�����	���X��A�my���,�f��EX����+�y�0�����S�B�_P����B']_��jϿ����#s/4[+��S�H�&��p&q��<#�%�;�����{�>	x���(���Δ���bAZ��պ��y;�W�$u��IኧI�N�������&[����{eͶ���q���M���N�\��{-(�L�1�b�i�펧���?<<j/{ɋ=A ��b^�������9J��^�g+�@c@"W)Ÿ��̔{Jp�7W� �9o�ĺ���q��Ɏ�_��������j�@�}����y�V�:d�@�w���BD
,|Y<
���O�X�T����,#B�-�������Q;z���;�E,�V3α)�FƖ�l�aC���A��#�U��֏Z��+g�4�X�??�@6�|^�b?�-A.�T�\�Y��LBL�.���\��#!�znj|�"2e�nR�+��\%����ϊHB_�A�H��o	���ы����(��*�!~bg�Nn�ׯ3:����J��/IC�&	e�-`.>����{)/����o�)����Z�B�����C«�d6q^���`z&�D�.�
G�NJM�a^��V�z�s���a��lnf�s����䐞��[6�Үw>���g�
8Oɔ��o�s��L��=�g؋^�b{�[���.�w���5���ZԞQЛ�B�əY?���k���$��Q��r�a�}�p��Y�7�Yz���P��*@���ew�U�r�j�`�\*n��_�����S�G��6��Y��cA�o	Yy(8����`�B�~�{�ч�e0����Y�B��g��{��y�a���K���w=#������x��k .Y^�Aۮs�p�'ON���H�јuET(�l�ju �{�s�*�X���l����`���BX,�
�!��Ț!HŻ�e0J����}�;((6��Ș����ȣG�g��M��S��>�h���e������ �v>����j�=�� �)z�(ޗ!�w9���k���0T`W0�`��������e M��DU8���9��;#��s��/���ۻ�ֆ�T��D�c�i�P�C��p��GF�TfAn����3J���V��@,�����n���Ea���Zv�����M�=�r������}ͮw�r��(��|o�˷9��1Q�P�P�� /�����(C��L�FO(���O:/��7���8
��# �Y�G���|���E1{	:���3��H�8G{�v�0$(����Lx#t�կr��a�V9��Lh�Ć��sa��'�&lU֭�>YK��L)�rs, �@�.)�i�2��j����@�.��V�;l��I���]1��`�ݒ�x��>+@�L���K.��5(���ov�"�2H�)��9�k+%S|/d�|�w=��X7��ʓ�(�����$%��$0xj��UK��%?�E�%@�(YJl.��$��&'<o�2!���,|^�:���%e �;�Y�E��?�"��^�qI]�>�*��<H�Խ��|��� �h,t�di�����}�(��	]�&�&����1��{��E�0_�����U����K+Wr1���mr_�kN3�� �'*ϰV�\�$�/������^h��2������9gqu�C���(���LLĊhkG�\����K�-˖۝/{�C��aR��c]��e[�f��ر�>����������A�]��ȓg���7�ǣ�x��٫^���za�fc�EK~ �~tt�Ɨ��-�0�*h)��1ɒa����E"�EJ0T<X�l`�}ua�9=.���W�,�bݩ��S,�4����\}*K�+�5C;�6��aS�ؘ󕅧�m��s��J[��2�2��AKZ%�A��M�~�(ā��E`Rp%:,Yb(A,"�K�'J!M@�cq.�T�у���TL�� �Q�(-�[j.�0`ŒWz(���Qr=	�r�Xn;�����,f��=�؍�B1�bD0���W�<�j�@��z�����
e�\"�	�4՘!�ε��P�j�.��X�֋��GZ4���j�Y����/��/�ڱ����x���;�d��������f��1���Pg��;'�,�P
JmOi6��4��i�}�I�+*��h�N۝�M5:��S�s}���� 2SN�Y�O�Ӏ��oϞ��>f�)���W����ړ�K�-�hX�ϸ�&�pi�hjjjL*/,c��j��9�U�8���)oϪ��Of���!�E�f�*�>Y�j�����{Ͻ���v�����Y	s%<��o����&o�c�E�1�"����&��g�gsܛ�A
".$.6��Rz�F��U���r��E]O#]�|u��5fO:��C>�*yJ�Sp׶P�Խ��W!��(�兒�|���UW�k���9#�j,N&V1����w�6%��M"J�h=E�%��EѢ8�.
��x��PЏ���pN	p6$B%�����h��$� ��s�������>���{'��MLsn��(R>U��w�f��1�dF�b�z?�M��:@��ޑ�z���2\R�����Q TEE��S�Y���KR�1��3KV�iv�Y�C�K��7J�NuY�:��KMg0�����H�����'ҘA�{�&&�����%S��$��
{�ہ�o���.'W�+|��J���
t�{�A��zXC����x���opo�����"��P��g�S�K���v��kS����#�/���o�kxN9Lz�u�������{1zX���G2���n��}��;ۇ����A�_v��v��O3x�[A�۳���_m��a۸�r�T���%���gϼ�v��W��@`�R8��J��(��Y lr�����l����-�4�s��-($kl��m�z�f��>n���¼���:O��w=��sY������a(���a�b�"���" �0X�@���{jW�k�@�3 -�{�E� ĺ>�7�e���`�J�?c�ca�T�~���Y���&eǨ��������� #��|�NA+\�j�9�h�sǺOy]t�P�<s ��84\B^V"
����?��� ���	�WN����ZZ���k�Z�>(k��9?���Ȩ��f1��S�ǳz��_�`���ՙN1
]�e/��4;Ią�����1�`���}���U[j��>Z���(���6ۚ���_a����C#nu:��V�I�����E��� ��w|��W�Ws
�=q��N[�ض��v�׾���
�t]�+"�i�БÏ����{�9w|��_����M7�b��~�ב`�T������/�����ٺ����M=����o�@�����8h�.wpjj�N��6�χ>�A�x�� A��sYQ�Q����	k���X�i%c�٢�z���b� ��Ҵ�e�e�k�7��2�x��0��sb���u��ӿ���֪Rf����Y����9?�!�U�L,{�9���_��s�4V5�� �ʔ��ō%����gs!D(�����a�X��<���]'X����y!��c�i����!��(&��uE�9�r�y�¶96�F��>����R��+HY7�(�aH�������7bJ��!�eaQ2�0Pe�}�e��:���a�k6����&\��;����2���dw���\�,y"��bAٙ�Ӫ�Փ^
���\;�|ݰ��s-��+�A��|{��[-��kT�chx�"kUƑ�Rd݋J�xz~$LM�8a�����o���p)��:�@��������W�x�����pҳ�%���i�w#�Y����T��˯��Ղ=���v�U��E�օM��Iϝ7?��u}:��e;����?�^���������\$d��ԉ��#�x�q�Aq�����¢��y�>z$w����}��[KV*EXyzZ1rxƍ���Ѕ3������rJGeQSEK�
x��d�ј�t��",��jD@#0�,BP]�Ԏ+�{�o6B��`�# �Q	�b)��S?�S���"WC!a�� Q��&���?ޘ�����X|�g̃2�k!��5���� ���>q� "`%�2c�\�ϱ��|��5A#d�p���)��Y��SS��+�eq�1�Tx:�JMv7/��%��En��o��1x�z�|�9I!�90g>#8�g�{|�S��g\����B���9e�Ⱥ��`<��G!YۋX=S�G���Z�زѱX���oY�V��`q#�wQ�ԝa���>��v������*������/��/�JC�!�x�x��`կ�fk¦�&���.yOP���<�^��o���*a��\����zљX���^����?4<�س;�s��:d�`={�CC1`Y���Z)z��MDe=��c�n8�?�s?�.?��B���~��XlJӫs:�?��n����O�KZ�d����U31y���3J�
�T%��$��9"�����H&����c(e���0 ���AEW|Ndp|����P 
�i��5`�r<��#�M-�2��=W�.�����w�����( )60J���#^�Uv�@H�(M�8�l�(�h="�Sȱz�S�[�4z�tXk�����=I�r/�)�9�p�0#J� �o��o��������yQ<�Ng��k����_��1GY�o{����\?�Hyf��{�r�5xq�K0���<	�`�s���y�y�]�(1=9�$
��cC�A@�O�G�@Φ�A9�xm@ ����܌�{NOO���
+Vm��q�dDF1#O�n+#v�gdU�&����1o���|��Wݐ�6�}�q�;d{v�
��B��jՠ���(�:k����{����r�3=^�^�:�}�b8Od����zc�1�]8��kqC� ��ix�O'X+v<ȄU_�2UySS'�����0p<��(����TH� p�����1�(-.�⧥�5�_D@O���ܢ'C���R�Y<cˣjV�> �P�i��;q���o橬���4�F�^}��2E8���%�l�3���6m�����íJQ-fq��`�����)}!��CmJa����b��+���ڎg�}q�W��ann&ǳ!��ξ[�J�;,L�x����q�V$�	]�=�ɿ�ï���9��������y�A���=�;�U�R�+k5-��9���y"��b�f�i�0w<�>���|�Z��
k��Z�
n�[����0��۰�yF#c'�@��ŋ뱩{��J 7�2���pY���`y _w�e����ed)u��g4X��@�4O�si��SB��g��r���}7<����~-v��n��
�X�[���!k7c~8<�Q`�S6��i�k�"��[��X�0KY�(�#p:0oa����h�BL@D��|���\�N��"���`���	�F��h6�R��4��[:��7�*V��)+9�#��kVPQx����̊"A
D�CA��V�Q�@�nZѫ�p\�V�'������[]��-*�Z̬�
`���ôЌ����֐�"�b)l^�󋋲Ty�Z~�P�������R�(�9?����MF��5�y��&���-�����P�����Z�x)�/J઒5-@C��$kIy���=�	����ow8�,1�jyF2���b(Z��w�M�ܵ���}�㠪�j�Ra��,8�?���G�v�X��Gl��N��iv3�:ˈ��N砤����l6x.@�p�?Yh��T��5�����+�jPp혵�=�v�Ѻ��1�Í��P��r�Ki�)�G/��y��!��y���d����A���j<�bL�D�V��)
5���c�P�	$�xpP
��	:;�!qq	b��>��M�⽲p�������c;�՜
�aN���i`�x;�zv���]xͲ&�=�(�S��`u;'��~	�Џ,e�H��yT ���:�\|5�Q��
�Dɠ@eJ��V�J���_/�%��*���)%�YB[��g�yu:?�PE����=�L�e��6���C�{!������ҌyaĚ�b�I����Q�T=�Y�7��ҕE�̓��	?��c����x�<��=R��A��ʘ�:ԁ}����K���"����}V��<�F�!�9� ��e��8Vu����X��O���m�v�� �n��w�\�Gcü���±�v���/5�W}�x��5���� ���(v+�2��ky�������v�8����������)���[zo�¿'m�,@��b��kæ>f�\|�ՃU276aa�jU�
�j��D����h�pW5��R�X,l򾱪�_���zVi�X��nq��M!���`��)=�}��F9�@m�f&OXi .��/D��Sh��螮�E��@#���|QG�k�*S�*�,��զ�q*�9����ɛ,e��m��;�D������"v���)��M+��{A*���'˞���NQ�oR����b���GE��x_�E�:X/BP�|GN�R'SG�S�'�R�j1NDy��!6J֯��xMp�FZI���EV����hR7�Eʇ���}5�)��ސ��Q
�7<%��p]��ĝ�_ۧ[���Y��X��	����7u��k)V���O>Go\�)�궜W+�Y���;_~��Q�"xU2��A�P��z����X�p�I�8yȦf��h<{otl�O�ѵ�[���=��9���h ���@����R���/��pn�G�n���%��+�28d;.}��~t��{�q�/�ff	tl,l�Ma��p�[�v�?��Nz[F���f�0�ʀß�?15i>������ٙ\�a�PQ.4��m"��o|�]WT�2�,�Y�p.Ulr�aA&��ȐMM#`��מ�b�i�}1�SV�E�()V'㪱{,,Zܩ[.8F�E��+�@l��(�=J3��L��������"}F�KiR�Bp�vJ��ІO��H	�t^��8H�C
�A�Y-R0e����|�@�E��\1�w�	
c�W�R���~��`������`�y���2�39硃G쑇w�.���*e{�?~�cSk���H�կD�Gw���"{��̯����mϣ��z���|�n?)��������>�1���
�5V������e�:�������O�/,:�w@>��OL7��)�mv�m��T-�{�1��I;r��a����t�^�5��K-���$7zPTp���C�R经��e�����=�����<[�9���m�}K_�re��d�uY�-7�Ɩ�&���m������&�����1[j�K9��˟�\$C�v�؃>ܫ�A��-��ԜW��߻/X���۾u�W���;qrʭ%pU Ua]���X�XTy�)���"J3:XLT�����qZi�܂�:2��`�dn}7X1mk461�p� ()�V\�7����J����к�BM��x�J�����R:x���/O3�FA��6+E(+���N{3��oY��W^�g_��)�df���*�:��C�Ǩb7e�1��
 ާr�c��CV��`-f<[ɕg�6�
�Յ���k��u?~�F�3�{ ���Η���V��}�/�ۺ�B�Fl��v�ȉȔ�U�
B\�v���b�����dT�Ѷz�ӥ�LƐ|����>�����F�e��I����^���UNi;kW<�Z_fG�ǵ�v���~�F���9�m�sX4XV�?�a����A��X_4W%��q�I{##hn&�2�����߽�A�������
��@���:	�em,�����^�:aِ���??��C^��7�´]tA��k�� �`�S�@l	�
�C��7��qA���H���(�B�ě���<(�{��R��|d8(� ؏��a���SRb>Jc�����?��n��\8�(�J�U,E����<�y�.���LA�³�÷�>���r*���&�0��۶^l/���Ju�9���q!��Zf#m�?�On�(���`�K�*V��T����v�R�g|��mlt�6l����똚8�{��ͷ\���ꫮ���"�C�'���͹3b�\j��¿k}�8*�&����{��?������k~��ʾ�m��w\7`��G����#I�t�����
���l��A,86A$gY,-|DiZ.k�J��yN�<<6��I���U���������d=kA	�J��XP�Ƿn��XZ�J��uKД�F ��k��De�G, /��18<�4&R��_�k��)�f1l��L 7͒b�Aq�7���]r��8��ķ����e�(��Q�U��K�}%�Pu 1!Ȩ�`�/:<K/��m[!^�f$�9d�ʒ�1��_���;�3]��& �Eߨ��}�?�Ǐ����g��Ipu)��`OWka�+3G�nt��k��=����l�5�7��-+�ݬ{.�<>OL��ۯ�{������Ïtء����=g;y������I�G�9�!;v�����ĭ(.鞠/��%C�u�����ұJ6��4��[�5�UF*x+/X�,�i��a(ȉ%��R
�-����*2�_�5kW�f&X)��
��9�aSԃ��n�*�����Tc7�蚗=��������4&� �A�PP��5(jkՙ`m�D��&댵�\�X�.��F��J�e}��N�=�¿�c���0K$�TZ#�t�K�{Zl��S\p^uv����d�n5�Q�r�@��g�'K�Y�1̼�pMk���.��r�`���Vm�ӵe�c����50�}�@'=/�����S��?�u.1>��G��j��P�4sQ��I��f� >���ڱ#��Ѓ��[c��68�6"�Yg������{����X���=����Y/��^��0{��ĉS���7�Nǃٺu�kjR�H�"O��*�͡^���ȌtNh�y��M#r~�|Xboy�[���H�� �U��1���
k��M�)<�x|��a�u��bFbN I��,�X�|~|���.@�X���0������ e@!$ș'��
�2߅v +{.��9>� ���M9\T_����W�@V�����C���J�5-�c@l((�c�߷϶���^�ĩ���^��AI�'�
H12*��^ĐY�V�����=�����͆�K�[τx=x�����F�!�c�p�����s��/X�6OTP]C��J�#����z��:�@���l٘�L����p�=�e���C�r�������l'�~E^1x��ȐkV�W�?��a�~���9�m�k9g?��MF&@ڶN�����]'+@�N,!�m���)�,k��+ћ8�ųe�6�eu(��G���7i����N�5�_*���`�Ȳmx����J/L�۰�y~�|e�Ɉm�u�Ќ�M��^N��6��5mө5�{� A^�q�7�<^���C�����\����<&�@��7�f� ��@)��0g�S�
���O�U��b���=�sq�*�3{�{1���"ݼ���k�>lr[��0s�T����g�Ůt1[�*�B�p�{�3���&v"��稩�~p���磔g�~�����>�E�r0�����h�2yj��aϊ|p`8��`?�8<��
�sS���Mr�dYɺa�@[1�փ���j���E�r�������1��Qx��%� iǔ�*��HpG�l��6���w�c{}�S0�cp�K�c;�J&L:9���4����k��a��!V�z�:�8���EN�ų�b��HM��5�����Kҁ��-9�T���lԱ����w��e�h�^_�җz���80�x�"���5��]�g
Ͳ�T�+Д���u�*�4�3����C���H�lWk��y�[�nS��P��b�K��xz�Vu��<n���*�p��u���T:��xN�� �r�ʼ�T���^�y�{�{�.�(��^�w�N�)^)|�Yz ���P'��[���%#�F�sb&-�/fe�N�fy�_�b(o�EΆ�J�5p~�a��}U*8'�PV���uc.|�+5��+�A[�b�M�<n3��
�����T��F����ٯ���K�D8 �`�KR����T ȿE�&����`����վ��3��,��CL@5(	������{�;�5���u�`�°��\`�:7�Tf�F��\�I�~+�o��H��b�9{�A�_�i��[���!�2�T�����#�S/GM
�R�c���m�2h'��AM�u�����}�7�tP��*�3��ꭺ����n�"M&sJɤ���(�L�������}V�>ޅ��� o��B�4�Rʷ��B�"��&�%�M��w�����:�H���q&&��Z
Mͳ�x���݂c��^��ѷ3�g�V�^^�Ƿr�/Y���
_�W�g��r��_�,�aQD �U�+�Y���`}i
�x�u���f�ȏ��.<Y2�87q+���y>G�&s��L�}Z����������x-�̤>~�K�8���ڧ��e���]�:Ԥ�R(+A��	�P
���v�N�H!�L��lN�c�O��{:7= D�!�������E�O���7��_8�D����WK6O��0����yZ}��7��]b8S��X@,l�XNlB�(cH�/�>�g�8�ڝ�X���d��˙k�ͨ4��Ջ�Ƿ|�x1��@(L��Z-�9.�X΂!����W��pf	
�S,��ǎ�m����>���ń��k�����W�5}z�}�Mp��H��~��6^A ��@U��b�]�X��&p>C!��Q'/)��A,�Ua�|�T�(/��N%bX7p;�X��r�t��WD*Z�V��ͨ�ݓ�#6T�g�gڍ�^,+R�g�z��ݷ�H���߽UZּ%�P����t�z�_xB����|"i�����v��t*	_̕�,
����S�8��#v�P,D#�'6���I2O<�y
�,��<��m=�U#��ֿX31��h� B@�����x"|�|��e�� %��Y�+_��(��k�@���Y�{<a��+6!��6�|��VsQ@$�b�s.���!
׈��us}�n�����Ҍs��-K;3��GOZ������И՛���NKy�q_f��ќ��p$U���PBJWr�C��!�o��}��3K|���z�U\Z����Xe����HcbStr��f@���g����]�}�6[�SCT�5��>u�U1����6�)n�~�Db=G�f����0����!�	��u�]��?��?��yV[f��8�)�|:r���g�������:��Fŋ�,9��S`]#�	�-N@��MQbc哵�<$������ �`�������z!c;B�Nk{���hp�?�����;.��1}����=�R�
̺1�윘f��+���b�ǐ�#��Wa1͢��su��q?g����ȫi{č�ajh�*�Gd`��Pڨ�r^�q�[/\3X�O�ɩ��lLY�B5�y&C'�T�f�K����dXv���v�����������3��e�,TQ!���:R� �bS*R���pLΑz��-b7Q���[�kJ{�w�J��G����`G��Ҥŭ��BOEe =~�u��.�0�V'B�@si6;�6u����e60X�L��R����S��~�=��RA�������k�57bY�w�l�'����	�?װ���,��h����قֆ]�*%��!KFCʡ�i�����ڀ9�s�C�Ϯ/^���<�Y]7?f�0�Ώo�L	Q`���N����4ax|�C#ܜ����E�	^��#G���NT��GP7�L9.1+�C1CF|_�\���W���wߝ[�@TdqM�3S9�������A�F�+H=Uj��STM�E��t%��Ub_��`FE^�j^��ʱ~Wῢ_o�K������HcnE'Xd.�ã63W咳��ߙ�H�j��ɫ����N>�؇� Lɍ�?U��-��ۨp��[��0SL^V:̅w��OG��H����O�)O�,����}Ѻk�x� �
�B���Y�D�um�`�5\Ѵ��ULS��� �v���S��Vp$�oz�0���9�$2|=�,�_���9�r*X�_�S����y��A>�&�K �}@�Z�~�&c���d��yۮGq�PO`�� HU%��'q��a���"�H��b��z� �S:���ؗ�={zF2rZ�R?|���޵?Ҡt#����%��2`'NM؇>�1�[+q�r)ҳ��xj70�HNq���8�����kg2�S�]�W�-�ʧOg�*F�`۳^�zV���ز����L�X���l�b�\�X��Y�~]�y&n��CG\H�2m�~�r�����Gg��I�+���f+V(f����>� �o�^8ǅ��Ӷ�SǬ7PX0��N=��<}�X-x�j^㪻���ȩr{�4�$��M�et]�0�|��G�A������w<'�Y��H���� 8��n�B�N˶|�����/��҃8�T��� hUg�⫵���	��ˮ
U�9E^E���[n����҅#��������Kw,踆��ګ���^��<�)pn?CŇ��87^FJO�2>�q�t#́��S�/�#|�68j�����ÐPQ��������V'�g�M��Zu`>�P�j+8w��}�R/8�\��G%�u�!���2��G<@�j�1[Y<�kE)׃bf���E6��l�+J��7��g��/�������lm�-8�7�!�O��v�~}�T(	��8(���]Ps��AҎR�"�Ry�ί�"�Bvn��e���v�ѱ����63q�]ڊpڠ�����v��1�7Z��o!.��OC�~��2t}*����L�I$����jCҴ]�wޙ	^X��)e�T�3p����%Av��AoX���sX�@5�a�"`��w�ݟ�����?T��^���G��H��X�R��<� U ��Dv��Ӵh-�����xq����+����Z9�^.e��ю�9/�(��p��XYO��� F�������U�G��������>+���Ӿ@�(�;�V���W\��Ä�����{<��޻��yH�����Ԟ��:��'�Q�S�*�p�c��\�dd�^������	њ��K����6�zԖ���۷�'?���O�J�E�+���,���jv&�h�������~�� F��ќsvy�x���#v|�DX(4np��J����-"aQ�pN8��eC�Ñ�/���,n�w~<�!.~�������� G=��D�),�!/(��5��Y���<DV���])"Y�b��wxM���f��*૶�i���֑��hX�Bܣ[�;y�n-�:�Pj�~�]s�e��m�;
�v���ܲek�˷#)�"B1#���6��R��ѭr�s��
��`+3Ii���]��ee�n��Y�������;^���	�j4Ȣ[�n�]{�u��ؾ��/�}��i���a�I���^�{D��۞�^�^Y\���ӮZ�?3;ִ=t؎�<�^��Uk���>P# �����0H��{���ܕ�7X��>��O{���:�&���`��Z��ێa,��R��������U�"�x'+Z���w� �W��I.�b"K-��z�<e�S���^N�x^��d�H����~��7k�կ~�c�<?�J��@a�b�s^�5�)PSz֥:�!�H�T�#�X ����Z���Utυ,.E@�F���9׀' ,�aD��9�3V��?�)�Mk�i�,CZ�Qw�(f����Ms���l�����٘v��z��s��@�o�{,��(OJ��w-S������x�N瀋��	o�>�Т�
^��V�U\�ƾ��_��_��m0����U�7sYr���z����.��U�9v�O�S'�z���������}�P 2<4jW^y��t�-62�<�Ղ=�Y��Ŋ++���@Ѝ�����@�
�Op�~}���h�z�С����o�ӥz�A�"��l�s��^���^@7���\�;��3�"DbKq?��lY{jB�TF��.E����xr��M��`�eRk{��g�D	M��q8���{�oe舁�2(�3����Ӆ;B
c��Y�<w�8�a�C���j_P�b�NF� �C���"@�F
�O<asF��c��I����7�r�l�!Q�_��p��o���N���Vl��Q+6P�ᆗU�
h��Uʶ�.{�*k�>�2��̝���E����a�L��=�;�p�a�^{������g�|����m;l����-ۂ2\m������c�֌�ٛg����Ӈ��z�_����ş?��˯�ʞq�Mv��^���G�O���/�q�gT�6�d'�����^��9��%�@)da��*'X�����������{(ɮ�\x�[�s����F3#�r@�H��g�c��f9��᷍��l�1^^��<�m9'EF9k�&O��t��|���s�ۧk���i�3u��=]U7�{Ύ��6�<����je���Mo���IY�Rs�̝�d͊3L�U��et�������?�	xu1Sis Kt����o���`�ca�} 3ȹBW�
�=?�%�aB_�(���H�Q�.J���C"B�j@��ר0� A�
���8����y��F
! ��~���8g2?���*��_+}q]8<R�EeP0`�1��4X�^�O�Z ��������Bޜ\���n��f�sޠB�O-�N#tC���4��L�RN8�@�2U7b8�f!N8-�\G�n�e���O�s�(;�C�w0�Z{ը&O=��<��C�k�.��^�z@
ټK#r�����]���x�,Y�'���Q�������cn<Щ/��z�����JcґO�����X���e|b�P4�5K�Y�bqT���?��O��x���C��&�Nc��R��8L��$�Fֱk��X��C�����=%�܀���C��<��~�;9�6�ɪ%G�`4�^,�-@lѕ�H�
g
v'�5���k������=7�	�P1���;`�d!a���I��*]��� ���� � X��
�TL��H����9�]<�&X�P$x���964�EL����E�Dx��H 7���Nd,�b�sa����f��`դ�W�y�j�G����Xo{:�^'}�+͍���l\�Z�5V����`�5,6�D5�>�A�HO�ׅ(����6��R�A��1��wE��j�T+#�����HWg�Tj�תқM�T�.G����?�o򋷾NV�� �V�4E�o߷�Y�/£�4������4�X2`M���әH|�ټI'z�2ٻ���.�0g� d�'&�TQDr�h�/49�%,X���〛qO,v4u�{���bs���l� �U�������\WW��s]R�M��A�KJ�c�D8�U�E
n��K�5
8�t� ���%*��%� �c��AE�nPldN`C7��P�q~���a�@���j@b�x6pg��W<8'�)�>1�sM�"�����H$*$|��̑����)�	�m�b�i�G^S��Ϫ�*�CU��Ra�,{x��}Kep`��������S*X��Bz#n����Z+Y̽\.�1\�=z�GO ����U��ɸn|�P�z�>���^�v�^GE&ը�zGw��G��d�X�cE�_��l���39s�F��{���q-�)/�-�6��BQ+�V�IOW�.��F��$��QT+n�Z����,��`��,-kzՄ!����P:q�:��Z�܍ՔH����w�i�6�&Zp�4'�[J�$"��jm*!��u����ez�hm�|,a��.X��Wb����,m5�^ ������sI�8�/x��$�&�V3>%�����B4�����}�vZ�Q�!��i���W,�����J�|�FXc^ ����������a(�C�^=6��v|� �C�^j��](��ߧ7�VZ��Ĥ|�d�����T��	|��޺�e+�������·�#�x1w0���IÍgxp�n��s�:�3���ۗx�&9
������y�]�s���M�����c�V�ϼ��Z�S_��3�< &���C����
�:�L6�`�@b�V�,Zj�<>�)��vx����}���l������©N[s��UX�P�\-
�x�FT�D0
x:���E��~*0�7��ix�e��!Y,~��7(YI�CқL�m�ϳ;��v p��b!+�ɷ��h,�:E��!Zm��S��}�����>R�gx\��a ���&�}( �����8��7�zQ��(�ώv��U%1X��~�a{���G 
��f�}	�j��`�խ�5�=��-�S�խiz�܂��
����rV��� k^@���?�cy�[�j�-6�G.�=(?��֮6��e8�
:�!
J.�1T!
��+�*Γ���Ge��{�
��x)����@��#)W���V���|.)�w�>��^�x`���QmG��.'����Q�X9ࡀ��ݿ�8���˧��8>��J"[�#��ȡ]r����EK��j��Er
��"RQ��"�T�z��p�� ��A����	D�A��ˎ�c���T���2�7x>��b<|�B����]�Uxn�,~"�$�'����r�}?Nx����Yx�n�v�f  �K����
}	��N!\#'z�8P>���:������nB����?C��D�W*��K��uOEe��2���C��t�%|����6�~$�VUϿZ	�=��S��;�}�{���pohbO����"e�'=8���f;���T���CϛM �$��>�1'�*�(F�FOθ�f1���9�S^��4s��ɴn�j��X��8��o&r\aUh��x�u]p��@�,����x��K�\p@䰘QJ�67-Y=����=\5i�8�o�^ߤdԺ��"g��8H�X}GӖ�v�K`���0g1�5v\�\�>�*?XC��;=dȇ������=IZ�P\|nx�a�@��eX��C�/��&(4d�� � ���%+������u�p�����Q�Qt�B�v֔�|w�}��
��q���ճ���o��8��)����Uu	t�E"jm�z_wv�˹[/�J��*�T���O��_�.)���@٤Ru?���½c�c[%naZ~���?�01o].�V��~	5��ať*R*oV�[#Se��Z/����i��~�m�w�AV7+~���~�*[�H���'�L�w�v�Ly)tvYy�Χ��2v��i�+҈��G������w�y���w��][����f� !� �a��tv�?2�o�BKf�4�Ua��EO��?��B\x8����Z����`����2QeT�~�C>�>�n��,ߘr�J�g���b�����Ig@4
�:�g�BKPX�;P�q����hL��a�T�����60M�F�9i�wS��EE �z&e�8�9���U'`1���H�m=2�����,�G  ȥ ��#���!�t�2Y�j��Ke5�ft�ܪ��7�vmM���5�\��A�H��}�z !^.��������X��v���-MUd��{e�sd|�\x����'d|�l�7����V������(H\��7�� ����E ��<������q`M����z�굌��ş�2z��1�4T�hp]�J.Hjűw�q�.o6\u�<|�zX�،p����I\��'6:��yv����ρ
�O��sD��B���0D����������v[�x�X,#�^*��|����W��(8*&�휺�p����w��@���>�)�V(BDØ�g�ٱږl��
���˩�V��=�#vC�����C���0%z(#B��q���l+a��6{`I�Ž!���G>��%�5p�}�c�R��m�](���P�ꀾ� �Ī�e�Y��[&�;�-�$j	�=���
��?�8����s���A6�K�bz?�C���iY�f����*��2tx���&&F�d,�.Hhn�z��u��$<?b�L�b��� ��͞������&]w, +��?�����~N]��y�.�$��8Ir��K�\i�yZCjX�ӷ1/�5�����p�c�(6g5j;����$.��a�ǯ�3���%a>O˟�B�,c�8�6"餱|��iE`�g
��(?���{���!A���Y?�����-�F/�`���U}�X=�%r�Tn�}p�O�Tq����L�#\w�QC�� �_��_J��0ҡ�$l֧� 4��u���Kj��a��AȝBΘ�׆36�5��h�ò����C�䓻��-���Fr�q���uq��>�e3/�FY��? _����u��U�rM]���iG<p׮r��ak�GͰ^��Ns)�q�C��p<��|�3�7�Ɋd �#�V�+^�
��W�l^+�i]�ӗO�v|R'��dCv=�CjU��֝��@>+�5���E-�T:�����Xp+�%��'(F�W�p�P���'��yQ��µ6����0"�Ճ9gXe����e2lCd�X��7C/[�Z�:��q|&*B;1��҇g�d-�E ���Bx#�okk�81i��By��l��R@�*Ž�F�#m\�į �݃Ec#�q���ڄd<�1�E:e׳~
4϶XQ��������A��0�BD(��Ї>��ϸ�gp�DZ]�{�!�6�����J]��d��@�����<8j�����l�v�z,��� %�m�}�d��5�i(x�q��V#p�bb�(����N)td�%/y��k9Ier�eW�Y��&IN6��*�U�����1w�?�c8tP����ֹ���k���H�R�����k������X��Q���]ۤ�_j�Ѓw�#�X*�:�gƅ��J@%�d�.�?�.�@�a�<����r���ܡ��pNl �5躓��վ�L����7��S����?���~׬Z]S�@y& Q�=6z̅�j�%䦳7ʅl3c�;`�j(�񊅐�� &�>rԎ�Y�0�rd�����{l=�
7(�8��EBki��a����V����P 𤡸 ��}�8�����Xƫ�Є�f��ի��[��FR>�����è��F�[^�R�3%5�r�K�������ռ�`<��/���y9�c�~�<����84��+��I.[-����\�(�~��!�c`rtJ>����C�<x\�x�(l���s�J���}�0�x0�L���p��T&�~��񉒹��t`�@�����pb�@� ɋ��x<,�~c��*!��.#,�|v&_���6���ŴI7hd! @��
S
�C���,,*�zc���D�c���  �ň\Y+`�!,�{D����m�/n�ه�an���<��>{H�;M�	�i�3��:,rҋ�w�e��_�m�ug�  q���7|���Hр�`]�<�'�>�{"�k�9(!��\ӣ���v`|8+W,�m�oAה��!�`�aF&U�wu�[���j7xwu0���$���ɸ�g쇛~��O~��	����J���M@�Q �	��,�[�J���$U,tv�cO<n��@A��!_0׋Aӝ��?��e؇}E��"��K�я~Ԅ?�
؜�dY��H� Ə���b3zǬ>,�?��?�ςW�f�|�4��bq�����gB��⛵:�B�T�'Tk	-��h�`Ψ�Q��m��CH���j���.�s/ ,0Z��� H�`�ạ�|b7Ɗ�����i|ZgZ�0&��� 7���7�O饢0	��[�����ǏkA��A��w�wm���_��	i6H��>��4��:X5�A�c���뿶�!��ϡ�PQ;T���&[�c���9���i�5b�sd^���p*�^�Z������\���s��z�"�^�|Y�|�]���S���j�Q����|����8��q����D����d��/����b��)/��d#$d.2�Ҙ`,>L>�U0�c��7,J��ȊȒo�ƳM#�}>�O��C�~��`�����;?��D]E��=$��b�r�@#�nD�"����C��Q5��mm9���h%B�����_h����{��d
d��j���XD^��/��`g)���>�|����h���a�\ ��{�]���a,����`������8'�C�<�������ll�C>�=7�R�,�FՅ�@��ϲ�{�T�޾���⹌�=��F	��� �R�*ܔz���?���9E�0����������=<G(W��^ �'�7�1�02�9������:��|�5~r��˰i�4�7��eec���Y���������0��I��k0�E�&�	�釞����EuH�<��s��0���Ca�L���U��2��m�ԋ��&|��ZG�o������m����Hos�~��o�+��aeb�A�����p,��/�.,�w��]	���!�������c���#$�Bˇz�ӦWɦG����i���<����M���Y=�U�@���7��ֿg���۴Y���K��[R���*�S���64�JK-UK���~��Y�HH�sG�������C���O����-���bIVi3�@�EzrW ��S^��7�Z�/Fg��������d�9��O���,6,�>�$P��d �Gr�%����o��L��:J�;��뒎�ZS�qݼ�p�k�}#���:�7��!��	��[�J ���Φ����>.��8�AC�\�X#C2n����7���a"EaϺV���%��3Ɍc5�c��B�'`�1@t�F�*����A�ǳR����'���w�Q��f?3�Dm�r��V�4�����m�:�+ӎ�>�0}d���������w[��Ph��½HXã�L���C��DC
���3f(��c���c��b�i/�1�L\{̰�9>���
�Ho��\�x�X�
��P ���U���[� V5?ϟ�l��l}���oTC)N�%�B��KnNʕI��fBG�4R�ؑ�ſӨ��F����n��D-�b!j��LaDWߧh�����rV���X}�(r�P �*��q\*,����J���P��	M�@������@1�G\��J��%��ҟ�]7Ce� <�??�R肇�ew��fA��y�汦,\j�9�_��P��q��=�1�"(?�opݸ�}�c���7�5��"�3�O���lY$��>�~=A+l�?N_��<��R�\Z�\d~۷Z���9c�<-��H�!��W.x,j|�)3�˦|�87,�Z�YS�	� ��e�?��q�wa'�L�l���j(�0� �AT!�,F�i9?l��>e,�n?&;�:k��(��!�?��}( h�0�DCk�	��6\��!b�T4P��nR�!1��3�l��ռG�Q��8��CD>�r����Hv�V���!��c�L�d��P8a���֫�7���q�?�9~��=����?��$J���L`ؓρ�<�$������<��fΆ������Nߘ�|�_�>'6�o��	�kCDxDJPX�'j  �a ���[@̵i�$�oq̮�&�՛����~�)�nE
9wO�c��6E��[D���,��FvōG+�����s��%�[t�3n���R{,l�����/���6��/0(�0����g���}�LBC�x��|H?��?�Z�~�����ѐ	F�/s]��ܵ.\�а��Z��n�\V�"0@�{F�����2�t�q�)��2K��h�^)ǐ�ؓͪ�E�\<Yw]4����	��g��)�i(����7&������':N{����;���VN�oՐۃ
�V�����	��l��e�p� I?"�=�S��Q� ��PO���ftb�^�D�T���F����9c���;�q2G�e��o�QPxFC̅w�1��\���;(MT�T��F���#�?$�HoϠ�^�A�U5�O(N��%��f��	z�T�����"bh�ъ��|N�"�@Z�E���IfB&9�,�ހ��i��!Z/P���s����T*�w�voeA7����r��n]��DTܗ���V��Cf�l����� �Q7��@7�Q6��+Z~�M{<W��kQ-q���ټL�F����K��ua�Fv���9cI^�74tHB$��h�3�O�"�3iT��4ʡ�-�8��a蘈?�C3ĕ��Ӝ�8��|��ӧn�`�#Q+��LK����f��|r�3yǇ��{<�}����ύ�$�,����T&[z�r�H9��(t��
c��b@Ӏ|�]}�cm��8�cv#��]����n���o88rW�Z:���V�e]]0ҜYŔ�4 %p�l���}�*x��"F߈�	^�b�:��̣�8i���"=�٨���4����  ޘ-.��Td8�w�h��°-v��|<.CA�|~a?��\�KK�_�R�ԪGb\+Y �b��Ѐ�Ti��LUʒ�,>ZE�_��u� �'���Ӷ���6f�I��v�t���)[S&4a�u>U�X�s���|Q[H��ܴ�vh��˷�����'8� �a�Ic�0�I �oȠtj�{��TP �L�_?Q�[��<O'2Ny�?''r<U���3���	.�����Xt�(�}aތv���Wr0���#�J�xD��k�f\%��
�TC,�+99U�kba������7Bc\�f��Ԙl&������h��5Z�HrhX�rprj�5H䆇G��Iވ���d�*Z.�^�W\_$v��'KR����d&�l͠��p�&�g�f�0����~Q��_X���F���?�8��f��%N�D
pChd�3�A�؊�������a�M<N
O�]��Dt��&u����bh)���D[��{��T,�F(�uߨ98_�~�]����I4��26Q�#G'��k��ϿVV�X�\/��M��'{�Ʊ1�T��w:�����ό�J��zcK]��K�O�I�Z3�P+�Z�
��:T�ҥY�'P�����U2Ĝ+:K��x���]�`}�^����V�Npq�fU��F�m˿����� T��1�6�\�p��er��73X��&�7M����y��կqpb��)Q�ҝcl��u�`Xv�6�Å!:ؔ��y����ʰD�8��1��;��T2k��U��C����%/�ŘH��5��7�~'�W�q<܁Mb���dE��>�d!�	��A�h��Ȯ��Lޗ��I1P�g�t�������6湟�;��u����毙�ol�56wMM�y�Ӵ���<���6&*����<�Y�ef/^����Le�4,z��Ҥ|���_��~/e��W�6?�/��[�o�Z1A福u?�@��1�f(�����8P��`�.�#�����d�gZ!�o�:����ϒ+.�\���oX%1��(�:����x�Є�iZ] ������U����'�z����1{9�r �=}�d`�Y��=�׼V�{�L	�(+��u�Ԫ�U���#�
�Ը�FG��L�wMi�Fdx��f#2%e���;W�V��b���d�X��K�����G��^3���
�f:���2��%�Gk@@4*��<���(x;���T��3�!�V�7{���ǧ�f3�ڨV�,�0��,��V�..�!"q>���n�.m>%g^Ohg�3FH�7�����$��$�%J�e�&��I��H�V^q򨤲*X¼Y��;0��E�S.H�����y�����y�E�P�J�)r�/Z���@��@?�D=Bz@�`/�3�Z�l\n&�c�PF?�FG9mI}�&�׆�J@�����u��<Fz��?�����"_E�������Ƌ��c J�JY3p��L��z,E��V�?,GF�4b��.3�4�'��(X����Z���L[��D������7��g2Xc�$��|�͇tC	ԬaRl��=i^X3���X�˰k!�]������(��aPV6tx�>�d�R��R��Ȧ�Ζ�k�[�� ��ߡ1�N�E��E^QԂ��r�
\;����*��ꄏZ��O���k�����I���/�X�ٲU��XeM���j�`e� �h�fO,�׽�u��YD���ˇM��D��d�"����0b�ȬE�o�,��}��45i:������czh>��kL�h�!�'%&TL(�@d�d:�_u�?2��@������4Bm���7��u��b�/�G7r���w�h/��y����HP��JkB�}&��#'\U���&�èG@��g2ܚm4 �.���\�}P3u`-��}���~?��*��ç�-���	BrhP
�j�|̏��X�7l��Q�h��dVn΄P�2���Ϫ������ร�_��-�E�Е+_M�=�x��GT���8~E�F�u0.�鄷	^���GS�h�X�O+Q*��8�c��T��p����}g�/���(�}�1t�1�U����T'z0'&N����ȇE�?�}��(䬝㱣#*�'�|\�������q�9r�ŗ��3j����?޾=!������u:7po阡�I� [��u�\�|��pJr�H���%w��=����K�汪�h�����^����L}@Xl7�|�qsӊ�5 �>r�B�;���<����_�z����[,c�� oj�+����Mق���"I�b¬h4��E����&������|�=��A��t#����ZY��U�(̙�`a3��1��V]qI�zL��n8P��YG��7h՗a�=4�?	��x�e���sq3�,��~���5,����F�	�Oڊ�,~��±��	Ⱖ�جi"OƦ/tmQ���҈��A6gE;
�nK����������R��G�� U�j���5m�tʅ$Cԩ��~=����P�t��$���g�W�<AJ�����v���,O^#�a���$�3��E�Y�<f��;N83��0%Qz����Y�C���k�5FS�����@oP���������߃�����7!{�<!�|ر�I+P��p�9,O��>����] ��Ke͚U�8��'w<������I�)/�[�}�[M��<O7�9��f�c�%���[�˭��"F8:<l�����_Z���{�g�a���2��6l��.���P�o����Qs�����o���a���d%8O���>� ��:�ıZ`Q�*�'�N�B�gI�,�����QF�$�Z��W��I��.����P�V���<��*��n�JY��B��9"ׂ̡�G+�!�{� �Z��j2�|H�S�:�[��j}DJ�q��(�5e���;oT��Vc�!��]X�8_Ը�(;u�"�%�!�jჷV�U��KO�R����E�*m��N��`mG�0�9*�ָ�U^�q�:�*@Gꗊ��Gus#�l�r΀���V%�����U3�d�ff
�|>Ãa��-�Vፐ_:t�j�ٺ9NVV��6���
��e�u��ީVc~��ǯWFr-�����Y��>��"��L�����`���"��_��������@��=����j܌���!��I]�����3��(�՛�*���-�7��笁;d���0W��
~�S^�����q�s&��͛�ڄ���ʷ��e�ֳ�uk����	�6fdl|B����	�y�u�]g� x�Gy$�h�F̎�V�h,�p��2f�����2�(�}S*�U�,D"�j�J�B4�=I�f�E+{���M��5 �j:���F�4�.<�r���g�/��Jy��+׮P!1�B<vC�p^�:@���ty�*���q����խ���C~�
��� E{��321Z6�epi���,Q-���+��v=.���p�K�8�B;+K���a�H��UUL��0p���T,)it˝j�g����#�^�#�s�'���/�;������REcޢ�wthJ���άtvAY�1<�I��g6�#E}��[��u�ͥ��)�� ϰ&��f&k��,��nTu9z����O�9<t����N��~,������cR���r>��I{,�1`U}cF�k_l����8b.�Ǽ�����n�[ �B���z�{�k�;�������=�\�T����񈮑��Y�D��)kh?Uv��K��������;�'+V���/���m�'���>�ih�e�<兿��� ���U�;�Q�������q:\(&�l-�p��B�S-�1k�v�-��%�Nm�����	�^ U��݋�/��/��@7%߭$wG3�ۉ�f:�f��E��I�m�ΕMg�։�������*�.�_7�V��@U��C�F�;������b�'��R#�.�ۈ�#uRy+V{��G��w���뮽J��ҮQ7�5��Z�D�#�������wn����u�Y�e�:U&�di����*��>V�o�^��(ʍ�]%}��t�۰�W#���kBqa�'Z&Ǝɒ%r��W�v^ ���\�>�HY�ꍤ��Bjt����#�ߴ������*.T���W���[=� �8�s5>V�o|�G��^p��?�i�/��!��IC�c�׳����m�,W^u���Y�9���	�F��R1���}Xʓr��[d��:?u����[�}ʱ��7��GF�^���K����<��E�����0���V��O2|�B�������~�+v.th����Д �������#r9C�航���xTe�r�?��q:R��2/}�K���蓣:Gw��r�%W�~h�ʕ�������f$���k1Ny�ߒ�'r�-Xh��Uj�8p�ڿ�P��֩��::T"n��*�qO
ZZ"����H%
��;�y�?��/ؿ	�d���\�6�
�|/c�O3���#maX)(�)�&�,*��zք�6>Si | lr����VQ��ch��k��"��Q�o���@Za������MB�%��e�S1���ʢ�	ز*�@/���`��-��p�f�︡�
�M)XE����q��B!{p���Y�5w��]C e@��oOA����Gz�s"��a�,C�j��u�A��~�
���B��Tծ6�BөF$��6�8!�Qu�"2�IxO�������Kh�fG��(���e3h2��zQY��	bNcsGx����p�0����@	�z���Hf��q��b�q3RH���kD������F$�eMJ6������L( �u���
�9��!t!C�^�7 �@����/����jҮbxl|D��R}�i[��a��	�$��󙔮�kk�DgGo���:�q����o;�����Y��h��8D���ߑ�!>��x8��@1��o�����P2l���|/����Ic4[K��ɒd�ŵk�yF9�؂��'"5WSV6m(���+"6mEh%�w ��<F�v�C@�@�{�X]��Z��[,��>+��Q$�1��	,$N+�)��ͨ�"1�#�آ�N@:�G�a��į��\�ؘ�rQ�6*��UХ$��}�*$�E*v�Z�b�]U,���M�EU�����nT$V 4K����ҁU7!�S��͍����`���K��T�~�
�|���ME�Y�Q�nM|`������*�lƞc��C��)�C�-}h�':ȕJS�iK�?_���3H�\�F�"�i�0��.Yh{*c���ײ�D�I�;K�B'��b�'
}�A`�{�{����ޒ��?��^�*���lﳾ�͎X=��Z2��^!��kA-i�$���&��,��`^\�:��n�2��3P�Tͪ&�R)���>�.�	F��	���v+�5	:eCnQb��+-g%=<�^z������7-.�������/}�K���`˾���}�9Z:���9�9Z)��,�kp/q�˨��E��*��:W�Ѕ�`� �Ě���3b��#��Аad �g"V["^\6��x,���5�Q�)�@b��0F��s�H��0��$���g�TW��6��nө72U���В�����d�D���x��A�ϪL��.�	(�sʚ�l?D筼���E�(��'	q�!Y=^�����2錛�c*劕j��	{�~Y�5m	_�S�u��z�����\C)�)���=8�qEP�_#w�$�[�<s-�~�O��a�Cj��:m�P�r�����Fw�>!�Hp߰�Br�gfM��c�Ν������oΫ����q���8�RdH�l��F�*U5�
�NWcr``�<f����=.'�E?����?�@U`GgA�����Kz�j���V�[�{���Y#���L��DE��V����6����^ ,�������K��+���|�#����\@$��U�ܠz�6}͌��۳5��������B�)uOIU���`�Y*X�CG�&�!���F"��F�j9v���\�g �[�`�a�NQ֡�fE̽��N����D�����>��g��ʆH*������g����1�u�������]����%a������5�Vv���W��UG��r�p��BcYU�cG�z�D/�`�����16Z���^��;t�����|%e-���hk�3��8����
Wmj�Gz�X��$�#g)�JU+�����̑#Cv{� B38�SQ������U��l~�z-׀�9S^z�\u�T&&;,��/��B������wK?��Sjh��W�hG�L�2#'��ǖ�+����q��gn=�Ċ�0�^��D w��;��p��� ��?k�~���uk7ȡ�g���V�����n���~����I)�|��[^���zpL'ͫX�8�$�%aN��54я�s�v��7�+�-W_�y��{���.��]�K,|�u�u�M[Wv�aX�F�W낯�ӟ����P7�t���o���0�~s�"7�$�o��o���E鉺-� p���b���˖���:Y�|�)��v>)�?-S��%E��EY+r��`�2Y�~��%�?�^FT��ԣ���c,�L�
�^������;e��5�v��1cC>�o�ZS%#��d:,�X�5 �*��'�fQ-[�Tϻ֊���{Z���%�)�\R9C� {_l7��8,��@��߰BV�Z/�� ���'ǆ����,T�kjD����������2A�D歹�T �-Y�v>*��~R�"ٲ%�%U�L>�)� B�%�ӻB֯9[ϻN��1����U>�T����K>�ڂ�)���\��Ⱥ���Ы����?�C�ј���p���R4�����}:��e�ʵ����d����Ԩ	�P�	sVL('t��Pa?�B�]+T���9����^��\6{MHDW��؈��4k�DӍ��j�}�8��1�.��ϱc�~��_��_���E�@����Rٹ�aٷ��Շt��V+��;��e��~y��'u�����,�F��@~ͼQim�EQx��}��#
m��bR�㮻�˥_&�j�#q�~�9rdhL���'�ʭ�1n�p�W˦�ےb�{��\>Ұ����`�����|�k_��Sf��1��s5��q�-�GN|D�C=!6�I�Z�Thde�곥�g�
�N�9��aCڬ��#G��sm�����L�����9c�f�����W�궚
c��Cf����X��D��2��@ϹV֮ۨ�YH�3Ղ�{߯
V��%��q�����w��sW��X-����JU��U9��rŹ�, ��^��N���M�.TA![P�Vz�d�؈^g�u���oZYU+W�wْ�r��3�"�ϓ�*��� @�*F��Qv�O*g�w����z7���*A���;/��R�Z������Wb�@1V��~�w�Z�)Y��G�?'?�~�
"�ʺ�v�zC׬�?��/���v�U��4 1ͫE�~c�����x<nq��-8�A� }Fh�۷\�:{�z =�,;{d�*���wD�1m��P�5Pn4�T��I����ǯ�hQ+Xf���]�z�z���~�����Χ���5�y�����}�3 ��[���!� $���սT���(���W	dr��Tv��~�U��s�7�h�Ȱ
�$\dJ��1:s�Q�Mҭ��#�������E/ԍ���^)W\q�Z~=�l���[�����.6K�/~�f���H�7��|�r�ԧ>eP:|�w~�w���a[��,�&�n!h.6���.���A�U�ꆯ��4fbq�n������.��YQV�ZŹ��~��4\��b��,��IIO�r�n�ֈɺ ��(O��c!�jC�Z�pܜ�TEܻ_��B-�^�2��M�b�UƻU��ˤ����T������Wk+��2���:u�;:���c&�sªY��l�*1�x����kM�@L��V]�� ����4mJ�����0�TC�W��֯�"#c���ڛD�4��F̀M���):O%��"�*�^�R\����H�`���z�=�dD�j�58�ӈg;Σ�s��J��Y��jYv�K�=�d�>��S%QO�1�U�T�w}E.o��z���Md�h�=�R�3�@�!��3:��~���X�L�
�Azy��y��F��Ac���%�F��<�P"�x��<�b�WR��q��Ss�2,tp}϶��ׂ�IՀC�����?���z��PBr�礝��<~Ȋ׼���[��,]��y���}�?�Ò����r�5�ɖsϓ��X���>�_�)����e�����?j%�<��U�� G�O"����)/��Fc�V���kn0aE�Sk'�ﰅ`t�z� �	d�X�@�� �9T��;��~�#y���-+W��!@iU,􁲦�O�2>Y_��X��<��,�zF^���e_'�ͤU�Bh�^��
��7�u����׾c������j��q�*���U2e�6�I�KRQ����m��yz�nٳg�\r�r����E��`�U`���{���&J�Id�����˱�1y�^��?_�EQ�mJ��
�@�W��MDQά�~���^��]�����ea�[o�U�٣Ϸd��(*������yq��n9g�6����S;���[/���&Y�r�Z��l��.[c��)��`�U��7�\6o�P��|�;ߖ��k����s6� �2B2��&�`EYl��h�֨�c�paC��?���ۥ�җ�D��id�t�B����*r5j��]{�z]c��#����9�\ 7��")輢�"�Ϲϫ�����R]��.ٲ�K�~�K_�b��oy�іXD�i��_��z��]��D�r	�^Bk�C?�ӞY��î}&@�R ,�\�
}�pѡ�:��S����ȵE��>X`����@fpO���� Q���A��k��P���s�̳Αo�9�������iN��d�$w�u��w�vɫq�~�1��g�o��=MNy�H+Ӡ�����y)����|�2Zg�;� �����N��z��g�����.��� ��g�/$w�	�C�ŀ�x�Ï>��lC�a,Z�-��8��%��	�@����Y#֟c��� �DW�j9��F������r>2<)˗ʹ[/�u�W� ,��ZX�g���Q��t�jA����19phH��v�
��,TS�ؽ
�2b��4�,H��D5�9����e�X��.�B�ظV��}��rV��87��0��eЩ2��Uo�wTWJ�l��X��b �ƘP:��0|Y��2}�y��'Գ�+�ܢ�|�����Vv=�A�!��"Jg����S�6WeAP6��@t��X�X(-g�EC(�]w�t� -�>�J����BY��K�QŠ�H2#4�0�Td��U�۷B��T{r���?d��\v��5�B���<G�0���e��Y�"/G����[^�U6��Y�*�.�Y�8�"��!��ݳD�Z�z+Crtx��vδyH�a�#w���q�.V�������9�p�ؓd�D�Ίeˍ��!_|�W0 �
�0��rYX���W\j�H��;�����s��##���ʑo盦T��;t�M�1WP˜^��K�<�pp������Mem~��ߕG}��;V�Yia��jo�;'���wВ�۷ߗ^r{�!0v��8>��Z%0*{�0�)|�S�4�Pr瓆�ս�	o��<���j���f�	*#n�r	N��']B�^u�!�9���㐁�$2N]-�RmqC�����@,�6�Ej�Ud�h+��JĪw+�X!mU�)K�A0cn�F;²�LNLY���c��ڋ�W����jgü�[��l�f��A�r��>���9���}��҃Ŗ
�"oČ��Ɋ	U��1cNZ�8�\6o���*5�r&x�:�]�H#�� �',i��@11��h��C�P!]��˲���c�5㺪��X>��Ƚ�T� }�g4:6ay�FX����n(��Q���x��F07C��y��F�,�B��R��ks�deGGg�9|�L~(R��=:iV�Ɛ�(YL������>"�"�P��8�~�Ϳjt ���� �9�����Y�c�+�
|�+_��M�e��.Dɶ�!Tv�ܽ��ͷ�q��ۿ�h��ET*1P�1�ZgA�����.�
���"&��V t��
�q��׿f�<�:� �U����x����ZR�0��i�� Uox������k֭�߻ݒ>��� �/��/m��B�G�����E<F��b�%����͊�@�WtE7i��8��u��L�"���$q²��nk�ё�!�mxR;G�GIP���0�՚��;��B](	�x�{n}"ǜ�U�?.	Cᙕ�QRp���¸f�Op^��
N��������g�{�.�7N�ȑU�K7�y+�r��(�M�TP�������I�0ra���Ūa]���)?\c*��Z��t�
�i�hV��P˭jJ7g�s�X�*�1Q��-����F��rE]��F��%��I$K5tךN�cZr��A �2����m�y_4��i����Z��>L�r?��e@=�?~ߟ�
X7d�>�Ʒ�������>A`㻀h�3�l��`�=�z]�o4��5BX00-�{�-	�#g\�l�m�>�[��X��c�R?RO,k��uu��B��[�(�B��׿�����`0"��'4>ڴ�9��2��2�4����a���&�1�npΨ� 4��̊h#$R��>.�g2nz��������n.X_��������/����!��^ ��@k�����2I�)�K$�`(���>��D">����2τ���["�P�g�OX��ݜ�*DQҎtnn)Zˁ	m�1 �,����"b6�~^㣅���ʙ�U�m��3�<S>������ߟ�� ���>�9�� ���D�^Ƴd�ܽ#�����T8'�|8h���s��6��aʹˎ!�3��Ȋ���ݴX	�B> E]�Ї�w����躄M'pY��\W���~�17]�t�O{ܪ�Y84�No|&:_���{Z��k��5$>����54�H�s��b�3���b�}2�{籉�'j�J���G�h���量>�-��AZp&�G�b�mmb�B�`O=�>��>�k����}�'��Z�v�F�욟04��W's�s�<�,��:�+rv�x ��>�,9�0|zOT4Xg8����|��8�k>�|�M��40��P���zh�aa�+`����O��L�=Sc�{&i-S�(Y��s�P8aP���rS(���>-5�"�{���M���~��;�w)l}�#T���y|AO��S���Ӓ'j������ p��2!Tدi~�|^�5�3�p[H�p<�ab��B��ÿ���.�G>������yoD�  b���-/ �
^��,����Ƃ� ��c����hNFs,�����ɤ7�'�m�i�yc�Vڇ?�a����}�����͍�>������7�s���P��L!�6�/�}�I���'��Mkʷ�\«��"6Z��5҂Ǳ���hnxc��y_�ӛ�s$�Wz$ �W����d(�a)���򇉀�����2���sH͖�o����}�~Z$H�4?,⯋VU긎�DyF~�g���-'k�f��u�w��N^��#��yDU?��y��ו�W�>���4p���q����O�
�h�%��Z9=c��
[�M<<�������>p�xA�#�e�^ ��6|Z�'{���!����+Z0��Z}��D�-�wz�x�gU�|�<���r��js�z|���|___b�3�G�L�B��p���A9Vw����������\�����4�3ŵ���yzE�Z����q�B�
�G����g���O:8�4p0'�(j��Q���ż�Y��+Þ�������9�=��Z�4<V��6�ۉ@�hٙ���Xsq/��/f��_d�6`% �	�I<
��M�\�}ف*e
!*1ߺa��0U4� �.9|d(&�j�X�͞�h���	�5�����c�3���5�y����=2|Ԅ�/����A�{�@b_���{�6L76�o��:g���Ő_�`}߁�"�s�u�b뉰�ߙ��@@�Ч���5%Z����>�(]�������-,��c226*ݽ=��:p�����87���8�x�~���:������>�~�]Ιڢ�c��:��,����Q"�S��[��g�dz���a��k��c��h�y��j��Kn$n�<^�uIRaa�c0AI4r���'�]��� �}�In��7�Ip�����l$b����L�����hY�@K���b��ap�O~�3�r4�f�Oa���.U�B��U���3ă�
!��.`�Y�CagB ���x0����܎�s��)�}t�����ߏ�7���00�Al߾݊S�5@1c#oT��n�5����2����s�d3��*w>_*zz����yP���<=��Ѝ�Ȍ��}���h�Od������ډ��L�Ml��+�u˗��Ń��H��p6)�
y�)q^�8�no��	&?]|�~8p�\�/?�����8�މz&�p�΃��_&�y���jm��9?��G��������ix��G�c���Ƿ���l(��0�
��6p�L��a���OC�
��Nǟ+*Z�;<��;���i�%Iq�A�`��V�)�4�4jq_+6#Qb�"�/�3hm>�� h�Rc��e�_�ͮ��<%]=�I�̚�x�]Za�d`�b�۱�ߌ~���Lt"j��h��76b�� 
����Ď,��~T*�d���;�8���<zܒMq��k1��s�a�#���?b��0����%T�I &�zg耉A?�K���R�;3|�����{)��x�����G��|�|��W�6س� �ņ�Oy�?Ο�/^̔_p�lݺU�����gYSr��!������S;-�%��'>���F�{��x��]���+
�V{��s{�'�g��3�G�{m !g�
D��oȽ�w�}VD�y�o���>Aˬ�ʳٔL��I�?/<���u����љ�Ze������p�g�s�>tD���;��"y���70�1�D�0��dCD����G{�������ʬ{1���g�^�k�J��_h�a�Zy���#i�a`":1��׹�|����i���J!!iֿ8��/|�M8NWwG�Ks! s����@ׯ_/o}�[�c��ii�~���Cdh��t�~���¥����h��h=f#h$z��믗[n���	�@0�g��-[�X��Aw�u�) �*,��Ny�ߘ��
`jr�������w�g�nk��{�N�x�K�ʦ�g�E�\f��(�B�6@�|�I+��
������_~����G�h_}�7�Bb�l��h��6RG4ú적~�K^�dFz{�L^ �������ADa��A��W��UV=��������F���
9�A����W_)��21>"#��r�]w�~U H����DL�<!�<|�zc�o��Tڈ�n��K����J�/}�|�ߴn^����jU�h�N���NȘ��o��h���O�3��W�C���GOW����ܿG����㏘G��R(�#����\x��&Pdx���lE��n�8b���Qs����s�\t�����)�V�etx�H�\����4���l-�j�>����ɫo�o���E\(w�q�'&�T���_ϻ�
��G��*��l;�<y�������޹K����h
 Z��H kBҎ��Vc���^'g�`�͓B}�g��^�23�ц!�B7t���o�Ċ��Rq�%�ʚU��V-�qZ�����cCOKg�*ݝ���RW����DE���w��񆛭��ٛ6�k�<��&�|���*�����o5l�!̢�}��_�ݲ՚z䳁<p�vY��G�ذR���ɤ�Z�i�6���P�~\?[S�������ꪫl1��G��6$�B^�}�{���7�2'�3���e�k��h�>�0靣;���Y�- r0������mo3��=��h�CV`�W+E��أ*+�j .�]�G%�	\߈L��O��ب�i����++V�1�Б����,>�:=Q�S^���a1�C���ի�J�^5�s�S�f������J��Svr������ݵk��t�M�;�Z��v[R��&ޯx�+l� ��\>(P=ca���( j��o��x��3�>��C�7�7I#R����W~�W����}��=],����<��òn�2�~���J:$�=-wv����49w�6k�y�g��e+�����/����-�g�
_8K��T0�)�I�VD[ɻ�O�oe�֤�!�0m�ᒱ*Z�����xa1@�Ӫ���+��������ϟ�V�!IZ{�G{���
\둃��;o������9~�������x����qR�<�{X����+�FJDVƋS�C�\iX��{�Tt�=?�W���Vk�T�K�Z��c!!�S^�A넯�42�M���{�|�;�J�h۵�C[?�'����/ ����/[|n����>=�y�<�$vj'|O�A�.l�9��G���>��gL��;�A�S�oذ��;�������-~~X�4�l�֟�0D���dJ��L8ցj��EǏ���	�5�Ԩ���,j�'lT+K��2����ٙ��֟4���0N�0H'�Ux��ĉ=8Y�����q�Xxn"�?2��]w��C�����0��h��;��Qx���ַ�%��ޝ���T�-oy�y�0����]�ش�'��P�̎�!'��Xod�4ʖOѤ�#�$�I�����r#�N�"�(j͞��4Y���ʥK,�a��R�Eƪ�J�%�q�1�ή��d�>�B�%~H�X����������\>򑏘�G�7�����Ѭ�����sj��>�0�[����~������G�O������˭��j{�`ޛ6m�O}�S�؊�M�H���/�5�֫LI����AQ��v�9I�p�(t��XY�_�m۶%b<f�"?�0[×V�/�a���
�y"�Zk׬R/��}�<�G��0�U��/.�JoO��-H�|P?7 �]v��e�>7
���`����"����=��K��?�qz��m��>(H��=컀����{v�o���MX�$y�������ꔳ��,�G��ɤ�,��υf�����6m��v�BG���	
F�X�q��iKu��R���]x�
�,[�R�ղ<��ӪaG�qG��!眳M.�����I\.6r��~`߁���|�8����wZ���ɇ��}�p�c�N�ʎ��q���W�'���ty��"��$V~GRg�d�YB�0�o�1[���,77)����8?�/�ɉ�K�������y�1�_�2�JƻX�J��5*  ��P�����Hދ����-$}��o �?&79�lbC�z2T2��gHzs�}!�
��_��s0��k�:�iP�����y�@��-��y�_����~��,��<4�1j�������?o�j�$+d�X��{:dO'��U���Y��(%K���_n�Q�����]O���s�}��������XИp<������=G^�����1Y�t�\z�UF�p���Y��T���˖�%����bIg���m�<t1$k':>������ :,AI����ÇfsQ�Q��h�gjpsb�#?q�����E�M�E��^@;�/k�B+�\�>ԕ��A�4�����m�=(x�~c�R}�/R��^�7=�`ǿ��կ���ߟ��=_1P]s�5r�7&�W���3���]���j�H��e/7K���&,2�DA��%�B�G�߉ޢ^7�F"�}#ȓ�o�9i��+<���$i$�U�A�1^�\_��WY���0#�a��?���������{����<�B��������0���<�ɟ���gC �y���׿���{��{6Ǆ{�a"$���"S�c�y��j�wȗ�����K�AC�=��/|�K���_�x��s�]�?\,��2��Φ��*��k}�s��z�^t�ҥ���yW��e�^���JZ5m���9�Q���6&������-��A�nX��n m�o��o�{����I�+���bwl�Mr7�W����!�[C52�%����䴾[?e�9���6L�h8f�7+}�
A:��Z���(�sB/D?\}�����/]�tV�����ph�ؘ���&�9ر> ��}�I���JdO?l7�kn��|A�>�LY�r��3O�^j��W�=��q?I]26���
E%9�u���S��ӛx"~��38z�b�	;�[�͈���k��<P��MG���,������gϊ�J?,��`�����C�����dQ���k��mF���d��+L�A��=��a�!��q�Fy׻ޕFrmq� �eq����TM���׾��\W�<e�RД��)�G~L����q�d��F�q�� ZP�<ɚ���7�pú��߿�v��B]f͆�=�Ѓ��s�w���L���zF�����#�=jud�%���~�*&
'Z|X���o!�b���UNE ���R�c����p�v�s-~��
����ϰJ���ߧ�dώ!!�W�ӨI�~��' �q8�^�{���`������8Y�ʕ��?/�m������}�[��l����=��a/���'�}eϵOO�k�ϖ덞�=Syvqs���uB@c�RI`��'�y*1�}0�_��,��y�fS~��{;�{ts�X)[A����g��/�����i�珌o������RR���f\!&Ъ��/+V�2W�O,���a�����zUd������M��0�?�iq�9n�W������l's����xa��%c�rȑ��^�|���� ^�������}sh�֧��I5X�xQ�Q��q�p��S�u����a�ؼ����xp����1i_����5���=�䥳Ё��f��rQXO�+9j9�T*�sCh3:o���뇑�^D�P�B���g�Y*.��(� �<BZ���%�^�'~�i�|�s��yŋ���/s�}��)=ey���>ԓ��~����7��]?>��}$b��Pq5+J�#��a�֭r�X请�[�T�ܷ�LV��l��~y����D��Z�I6?�C�NS���rv�:��\�!~%� ���?����d`�	',V$��.C01���OǌX���f��}�!x�,xp����7[�>� ��O@���͍͌P�� �i����`��%�������7==)��5��7�,T
LB#���~7���$)^V^��ot|,��)@1�D#1�!6�zBPњ�9���0mV���9iı��1{:{���B�����Iٹ{�k�L�/|*&��=P�C��8��g�|�)��1��c68'�p��s�����g���3`�����b`?`��0�9�,{V��y=I���مD�yqo����tp���կ�#����~�~G����)-?�Ž�^޵F�x��\j �B�^1�a�����G��R�Щ�:���N��F����?h�v4n�u�k.�6`E�Ʉ.�ѝ�j����|GN��,X�VD�`#�DՇ?�����w��xӛ����̈́�/�N�`;J�#64��f�Xf��惫⸰��=P��l����D���a�;=\6�e2ˍ�����I,��}D��+�(�yh�IbZ��Vz/��1�ZR�^�C�E��XQ��h>��r��C��,P��J��*(N�p�<��,p*�f��?Wț�ea�8yJ�M����� �`��s�;��|��dqds��� ��1���i��� ���F>�=L�����[z>Jέ��TPիr���A�,�$k0N�Cr�5����ú�0/b����"	,�=91e�	���U���I���p�$q�t�I4�ߍ���X�e�2 ��dŊ���Й78ق���k?��w1|8'��ߩ�����r|�()X��_h�j�Э���q+�D���q|��6�����0�ޜ�W����(`}��l��Ij^+Xb-Y7�0�C\�)���{�� �,H��_=���{�Ռ�3gB��������[�:����\�0�G|v\���p�?>>C�|���S�g7/��J��珠��:#E�%�ߢՇ�b-�o �d2j,�l����&��8�,e�dB��ϲ���{b#h��u��ۨ���?V	�^d}1�0m�� �;Xh�]�X�hcc="��x�ܳ��f�=��C�@�x�Y� a�pQ�R���̑l~q/��(nf��Ru�h?��j�q�)���KH��Й�}V���%��;@ZY�R7��������˾��i��L濓�ϴ9tJ&�vt a������)<�P�<5�����o?gp`�#Wt��Xx�� �\g&��D0֜����3	�3p�����Hl�ÿ*?�M���8����l:cs��17��ʦ�4�e
�,��!�Ű�M|���,�<�߮/�p�=��a�{°�	�<�.����u��3���	�`��&��ǉ\�9|�;�� TuA�Z]zR���w��m�W�@�$��� 7��o�/}�K�w�ð���c0��_���>��ǥ�ǩ=�}�C��
a[`�ִ�o�qӷ��~��k4b���t�7�ik×ʹ�?�8兿�C�0s2�sq������`��ۿ�[��9����p��C�dl�H��!������g{L�F�
lME���j�z�=~�G��>L�'w�3LO���A�������� �+fr�
�f����9�F��D�I�8����6��)0��1<?��G��虑	����d����(L�g}�b�q���sz;�<��6�����Cs���������W���y��<������V$�O�q�8�HY�|O�3 Ny��A}<�`6������b?�O4F3���P���ΰ6B�D�l5���������`��,n��(\�h�}�͖}̤S��1�n�3n<s^�1��;!���Oo��'�s{�c��ii`�u����`}m��Ux'#r�ۢ�+��)�g.|���'�����M�4��h	�0�w��k�w�l��~� 
��
^
@=�io��s`���"�t��|@{�,��Ѭ����_���?}���Ж�-�F�	|�ٺjSP�{|�%ףUT(�ݻ�����B�R=�P����B|�,��9}�d��s�܍ފO[܌��B��z����MFG�J'��Dn�|�x^=(V�2\f?��̦������|�����x�,��I�XC�b~�c6�?9JGR�T+�����������r����>�oQ��lI�l�7\�1L��I~ ���Jȟ�E YR+!�$� �)�1`\0`\�1��]�,ٖUn�w���g��9����;�;��+m��\͜9�-��gW5�?���U+���bZfO�*`A�Ey����.1�l����[)��a�;�l�5�GaY���H(���cQ��p<�-���k��7����Y��{�ޅǰ�����"�{��P�4�y{^[�w�1~�����W� Vڣ�#�}c�+m���?��UuN�W��ZE*e�|Qq�^�-�w��m
c̊;l �����+�u'j����2y��؊S��Y�ąN�*�����8
��Mt?!c��D*d%�ez`�<m��1X� e��8�}[������0Xm��%K�m�p�Z���,��D�sT�����sl�$���.F�<�
���3�56Z��(bKgRzL�Z� ���#�(1p����JX�F�A!Bs��.P�Z�� � ����Fh�ز�N�b�(qL�R�1�B���9f%lR�v����G��9�t�b,��7���x�	���8�}.��sj���ϙ3[Fǆ��zp���A�]~��q��ߢ|�VK��!�дg�A�WD۱�0Y���}�\v��N���Z.)�b	Mݻ
�Ig����uN  �1 @�l��
^�fc!��Z��GX�YL��Iu�����&��N�Q4�U`0��Lm��u,d��dT 2A�q`�)Y�KfNm�V���"��Mgb�:��Η��,��d��r�S��N�	��1��2��Z"���ñ}�5�Ԃ9~�'��ٓ�<�!S�q*
y
��5Pج¦���R����� ����պyO[0�}��h�A�ь� pOj��5HAa�/�OXw���7�Y�
>��,=�9�u.���Y��sf͒׾�5���\���^a���S~6��4I�Ƅ`�g��`yL֟z���Ȭ�3�f������=�ec1\��c����9�Md�6ky���._���b$E��� �a���B�Z�&��D�$�؁��K����d5C
4ݘn��Y'c�8�#0�!5yj�d�8?z�W)Y�O��M�sw��59���ٳba���иy��[�%
�;�.BQg�g��92�����b�3\PL ��X`�cQ� r� b�>�bT���xˠ^-�������G�f"K�L������L�������a��D���&������cl�P"�Nz_�����t����]�O�tQ9!��U���_�����%�8��ݷ�٧䷿�[��t캻���h�)9��c��7��u��k~$/�� �@z��ml�i��C	�z�8y̓/<_�͟-��N����~%[�>+%'�!e+���9&O<&3,ǝx�t��ҎPhG�~lR�?��]�SN9E���_�m�K퉌����$���"2C0	t.BĶ\�ϟ�-�;p΁e4ٽS_�j�\v�eu�t&��Ʉ�&��ǀ fs�A-���.���Q�̟Z�O~z�jRV3�1�
�L�-'ў�`iDs%�0 ��o�a��Dc�p�b}��K���.���C(�X4����C��U���M
e��s�9G�=(ȒZ?^�=p��z��x���S�Źѥ�!a�R8[��>>��kY��f�{B;�3�<ӯ�Tz�rD`3��%q�/c�A��ޤq.4�w���O��|`\<Hm ~���uD�� @;̕+�;!^t��O6��<������(� �z��k�rB����M���;������B��`��� ��YS�  �A�-���\9�%R���}���e��s�;����-�����'w�u�l~�Ey�;߫Z��@�>9�(�t�^{��7����_�z�h�� ��_�<�7�abc�'�	'�0�1�Uc5i=4<S�����8���<�+
�]n�yO��غ	B�q�ʬ���jo��0�?���4��P�h�y�\U�����f�02+�0&`Rt���E{>�#�9s��r��hL���)v�^�����}�m��*��i|=���cM���E;�ItS]�c>)�gŊq۴�������Bj7#��&�׮�S�y��C��82ִ�]?6 ͽO��Z����ZQ{��1f����G�޾��o�J	��P��k�S �,�?z�<��S��9�;��~��<������ʍwEN[�T���=�|y���Um�|L{�6���is���渍}�G�s��;n�#W-��;�ir�ed�_��7�G�B�� �<ޠR��6���>L:�p`� &�@7h�hm���7�u ��6֯����t�n�6H���b�H�9��[_2!0o��Q���vM�ic�Wۀ4�),,tv�����b_./]td�60=Q6�2dtn��|]O���0%�źk+_p>WPE��@ 
��1j���0F��gLJ��͞�-3�5�y�:����S+�A�ҹ���x�Y2ѵ�?�k�
,�Mco�8�vp�úB������WW0�� ���|򓟔[n�E;�q��~a=�=��?%�g��Z(7=	�(�+ȩ�Y����W;
._v�
�#�X#����[;�)W�N{��,ϟ�L��×����twed�K/ʑ+�Ȍޜ̘�U(]��LAd�Z��c�ve��21��܅	�f4�|���Lr��.��b5��XsP+AýMt=�O�m8������l���7HR�M4�z
�����Z��q]��O����y-�O�I��P�4ux�
f��x2Qjy4�q��lf��d��k``� ��x-��6�)�`��ٜf8"�}#�$÷)�d�xv4Ɂ&��r���B�)����^���Q�̙׎!���ϛ�}p�����Mg���|�l�5쫽�?x~�g� pK�.U��������Ö���B�p(��7��`�6�>"�g�d���2w�wÏ�X�hA�����-ȝ��[/\!�3g����e�aK���Ti�3�f�����F��;G%l��-۶=�-HA;F�v�;I���[yL�|�8�S�`�Ϛ�AƑꈺ
�����_�1����Њ��翐����̙77�Y??Lln��I4��t�������y�|��Ǖ�=&���s�E���q`�b����:'s�)�d��]�
�����X��6��f3ڋᩧ���$�;�L��ܺZ@����70(���������3 ��
w�r���)�C!±��êD��fy��6&���঺t�z���?�-/k�P3��q��d����a�ARY�.*úRk���M�m��b>���*��C��MoR�/�� ı  ��s���^{񅗜U��?�(�g���NȎ��q�"�q�Y��ky����.�M�����_|�y�Vp����h�3�Qbb�v�ʦs��Ckԁ��lJ��ɡ��c�5�ӒqǏ�n���Q�ƄM�F�^2w6��d��M�l�9��=a�a<�,��5*���V����O�qܬ`�}um:� �^��8��Ա���}c������cj���6va��Y"w,	0�fy�,X��F�<��gצe����%ƿ'"��®++���I����"�f�q��ʰnЫ�3���|�󟏳�p����ަ�~�/��8]'N��#w!Z6VkN�G6W&���J��`�qp��)�t2���5�6':b<��O��B
d�8�ȫ^v�
��g^�Їv��wҵK���ag��iSK��;�ͬ�X��p饗j�j��@0��{�y�7d�gf�X_��$n4�dL����J܂�%6�f7>c��L���[�i}��\N �1�c5P�l=)sh���8�3�+��
U��-�i�67����%%�k����c��4c�v�9�|>S2Pm����#�wؾ���xnd���_��j��v���������g?��c|i�0#��B����3*�rF{���ު��yi�Q�@]�iY��-�Ҡ����S"kHR�0Г������x���	�_��	�/=��=g�̞��i�nӧ
jrժ6 ��K���\�Grd�5�ό�{�G}��}�k��;�6rva~�+_����7�f�Y�n�6���Zs���u�-cO.�F�d5�fZ0�ϑ<�-@%���Lx�d�Q+4��B�g5|^�~�8s�h�Xo2��˞�ײ��^׎�i(�~3�k����K�}����J���L�eb���e@7yO��ܛ�k��`V���뿎�'�� Ա�Y���cb�
�×.��b5-�l |"B5��I�`����󥧷�E�>�E�B��[+��q���?&o��5_������3ϐ�;v9F}���}��9)�#�fuG�+9YԻ��Ԟ�.+V���-$9Z5R+����P� r�!>����>�1�җ��ھ�ٸ� h�l�7�'%�o�_��%��̈́�ua�sY��M��Y��t3q��2jF�1w���|�y�6Va��V�?��y�ɿ��������
�f�׎5��H��9��[?=�����co�CA`c1��j���]�E��MaGK ��9���{����p�����@	��dՑ�ep�%���B�L�vVB��U�Y9��3���k6�G�@�>�X���$޳�0L��P�����\Z�{��.7��{�L5ǰ��966$4fϤ��v��r��r9�����0�M�6�@N�h,��.�*`��?���p̒a�������,m'�!��Z�e ����2U�:HZ�>�L�j��Ѫ�Ԉ�l�E���&�߼n+���&yV��3
C+x,��cb�Jj�,���P�ot�V,��{.�Z�1Ѽ�m���B���(vC��;3߬0~�ޠAw�&p,���:J��,;���T�Y�R)�M�1�h2�ͻs�e�;�s�tǮRK ���[�QQ�k��:o�WUZ��r��r�mw�+/8_F�Z�d���"�������c
]r�I���^"s�-t����wOp���_���wj��~�� @̶m�����l}���bd���w�/�9��i�$����ؤ�8Y�����h�[ �%��O���ǤO�5b����`�2+k�7Ҿ[y������3��cac��ڠ�T�2�F�9?�ț�[]TlƘe�������v-���������KZ�M�EV,y$s�uI%�{��塇�SO^'��,9��N����]���������b�r�y���k��r1����]�=*]��b�Dn����?�?I~� �'��?��P��c�s_����\�������ŭn�f���9��8�U��� ����=�,���0�9|���*�׮Q낛�n �q�O"^�D���Í�{�I�}���=�s翭��U��H�p�m�)���p{��>R��粩�I����
~N렙�k�u[��<&7�s�T�Ɉ�g�xr�W���Z���fa �?��?W�>g��f�� H��;{��\�J
�9��3�UGɖ�7��� %��L֬^�, �SR9�%��#���?�ŝ5.��s��V��=�oF~��9L��\u��w�Z��	��9G�Ξ[߬nB�ق���u�}/�������?��?>G�=��ƍ��͛b�.d���.Y읤o�L���`l�2�F ɸ,�� �����>P#�ОR��Z�7I�����ͮm�C��7���jF��1�&��~��o����a�k�m��k� �}?p�Dw�2��ـ�����A��
O�������7�M?��gH�[����I'�.���xP�]#x�P��n����:+�?��� ���S|�����^�.`g#0s�q�)�6�}L$.��6l�GyL�=�0���l,�w��ݺP�@��8��?��'�.�={v�;5�v��� �8#i�X�8��QV�>D��`%�ka��}ٲe��|�f=��E]$?���!�ҽ����{?��b;�q��b�
�'2��/bk
(N���=���Nhx��g*�B�z�N@���u�W� S�7C�vI��}� ���u� (��[�@ ��>@j 4���|�Wj��Ƣ @�> �z�ߨ��XP� Y'���
�/Ns���Q0j �vb�:�S�a�#U�C��Z�@�E��x�`�Ŷ��a�Ê��������C? �;aR�g�2�*j�V��R�r�_����ө��N�N���G0�Aq�"Xa���&
�
�Dj*�7Z�����& x!ЋB.��~�a�馛tB�����f! �:�����Ad�eQH�F������Ƈ��Ob�������ܢf�+����˿T�
�u���� �l����3}'����ξ�}o��4SWÈ��aӞ�7���<`pA, �xV2ٌ]@�����t2Ku@+[}���h�$����=����;��&�M[#=��"3�=D��`%��2�M��1����������` ,	��{M�E+�?���� �֮�����[��gS�q�FA:OL�g��|�8�!���Zq���.��-�3+�S6�[ڝe�������XT>@�"�EĎJ6ۢĸ�f��%����{��E~���v��!���p�0����}�s d3�\�f��dVF*^ڗ��BOlex�>�k����PZٞm�g3�OGn'���R� oZ{�z�|��K�4���E��v���_�O�ӊ� ��XLHE��׾��* �o���ЮۅZ?�6����l6������=n�OX��`05||��O�~��/����f��|�+V|L�1`��
�y�@N�{��LZ����'���D�i�	���g�M�����]��N@*=��"�Whְ�̜Z�L>�����҂�}���"J���4PJ�$FK�f~�h��)��ŋ��� �������E�<���5�O�8hNcކ��ֻ�Ѻk��`������ҩП����/�l���m	2��=��f�Y�E�3�#�^����7[�kB�q��>��<]�A��{K=B��/��h�	�+�@�J=��~�z*�׺�ƶRZ�D�02��@<V��oP� 0bҷ�ܡ�$ѯ�ģ�3���(��^s��=C�;�X��e�M|*���y�X���cŇ���@d�X��Np�=�j��e�,�T}+?x>�r����z�����β��J���촞,Vp0E��^)'L��3��� ���ZM��N� �k�]�ijn��1����� ���[�)����U�xR���@�琡ں�d�� (�$Pf�AV�K֊���bƎu��,�m��?����[z��]��]�"~�N��sLg�S�����L��aJ�����[�!�hzІES�g	�,w��ò� N��G�x�z�"��Mz�p��DGc�^K��s�0��շ�yj�48'�o�vl�
ٜf̔��fh�K�k��cJ�RHd��E�ð���;GB'�*��ҹ,L7񚿿�={G+Č�`�Kѽ�:�e�J9�-��0�}G�����/�K�_���71H��t+�Aºd&W���@!�%P���s����O�Ly<{e`�����R3EN[�"#d�5~>�,j�_���ղ��T�h%���󟴁�����5�)*W�:I�5`/GЭ�jݯO���:�m��V�"s�����M�DR����A����YRp�*�����O#�F�;����>;%i����;�̌��B�t���<t�8�T�u�A�,��|���쳲t�ar�y��9�,����NP k
̿
�B�1�ZQ��[u���-U�W���H:�J_��|Ӎ
ّΠ�O&������q½w�*�8>��F�,5��}E�_0[Z�!�M��(`�x�����T�|�[8��dd-�F�t+�L ���5x�*nQ�O�[�,�EJh���i��C	�b$@���ה�����3#n��H��V5���v�I?i^'K��6ɓ�k~x�Ө�ҋ����n0f��i/�]�E�Z��eo�_J��ݲ`�|��;�i@�R-"���4�XK2�Ǚ��;�4�Tg������E(�� ~��3�����	*���䶕���fc�nӹ�̘�#��,�o��Kp;���@�FF��B��2P$0~:P\=�p���&�L L�%���SH4�R?�J�e���GX�z���zu�R�F��z�(�<nw�Z��k�!Ϳ!�}zٰ�1�rMq�1��C�n�u�.����(���}n���wO]���mTQLַc�{Β�YrQ�?�}�i��%g�h�Ϩti�W�� ��,�h��~{�/��Iw���Ԫ���^ɧ�B�He~xǂk���!��.�9&0�"NVkS����g�?W-�� ��T:$�ZY��9uE�
y	�Z��Q�����"�XM�ʽ8U���Gx�LCf=�Ex%fՁ^����
�6k���Z]�&C�X��w�8X�*��4Ѱ��������5p��A�=4|,("+
����n��w�1�Ë��M�����	[���b2�}���G�9F̐l�G��Uefź�5W��xn��3��*B�^Vj�蕙s�h���`���%�<:be�7���9���gܳ�z�%ǐSmdD��i���ԱgYcN<S�FS���	�J�397�9't2��S�b���|�ΠӚc��D���0�FOk���`�׶4���E~�Sr�'�1��؈,�?_+���fb\��B�W����6�ӰKQK�\1�������>�h��[�MY�l(�)��ŗ�RN?�tQ=0J���>�9�u���jr{ٮD�dU��Pۣ���Į5.�ae����$К��������1�*�����o4����vz���hmX�8m>���T��y��s�Nh�Kge�1�.�}%�I&�չ��v	�4CrZߝ���
��sK�{�.'�rRvB�\)�X��!˖.�MO?�kb;4I�4����9�:P�%d�̘�#�'.�Ŝ�3ئ�:5�3β>��3��sϓ�n]A1�
�`~u��ZIL�������}M{���3hJ�ޞ�����sΕ׿�5Z�U.�jZ$�%�"r!k� Z��|��_��6m�tO[���i�j���+9F��c����qV����U  �"�;E��ct%�}���p#�qi�PkN�h��H���tI՜�VH���G�2V��ʘT���v�;�0�B��˘ȔR=5[��-Q�eU�⳺$����L*�Wh�1��~֢� 1,�c�����u2 69gS�|�Q��ýv �Dֿ�72Yy��ީ�������ݏ������w) ��UGʯ�k��m��|��.���D_L{���(f��)��"W��M�Q:��M�T�n���"}�}�`��Ys��Xy��dg�q����ۿ�[\-�I�$����?��?��~���'�&�ැ�>L՛����3L�Q����n仫pH��X�� ���{ѣM�8�B������$,�J�����R�8�;�>K�J-3&Eg%Hۚ��}G_�'�jydB��H�+�Vk("s>@�T�9�WM��+O�������5P��n�U{y�`2c��݊{���P�t��u��l�e�{��J{'��I��� ��Ś�~���mJ�e K�{�ʕ-��P�9�����K��a�ڬ?޳���1�������6Y�z� ]�/tV�}�<�ݼ0.,�#�X��u؍UY���Μ��f�k�<2�n�3��ɾ��x��*K�,��^y�t�s2sV�lټQ~�>y����o��Du��'�g��Qǜ �ן����e�]����s�9��կ�a�� ~�t��o�]���oi�7��Y"֠��h�M�{J��:t�F�J��8���0�i��U�V�-�·��L@�&�]x���>�.�2��Z �4�`Yw���G�1��%���R��ߖi��Z����tYw�M��.ٚ3�L�%�J>�M�`�<S-z&]BG��Y+�b�St"���H�<@� �
{�9�����p��_�=�0 �/��r9�5Z̈ڢMO>��Z��9�:�v�nY�r��~�ٲ�5�,��;Y1�  l��Tb�Ӟ�7#g89�c�`h����Ҷg���[��#����h��Ӣ�����V����}�yH=��3�_ߩ�`,
hӐ�-^"7�|�B�b°@������=��3yV�/j+,m�7�Oj&)��\��(�pZc>�6t5#���K���s�������ˏW&���VI;��7橥*�ʨ� ����^��� ��J�$�6��d۞��m�62(��j{�&�M�&���70��ɸ�M���?�LP��ReS[=K8�N=C������rꩧꞇ���/��b�����=�ZE�ݬ8��ի���O�տ�rܼ�Qyⱇ����+�?,�-c�J�������ΖSן�	
�7>����r��^'t!�)��g�M*|�Y��*U��a��淿��yY�l������^ �<�B�ᑊ�x��r�jY�x�Jx4kA��>K,��[��Yg����������?_@<�І����tM��{*�aG�Qq��|v�P���@Z�5rbld؍u��AT�&��K�?��?A2�j�pM�R�Z��u��b����1�q�5W��ـ!u��+�Ȃ'2���2:��0%�{��G�s[�oߩ�C�c�ȯ�JH�H���%3��;:�&�e1ЦA����*~��R;�1J�C|�d��?^>��O��c���Au����~m����^}�,�x�*�]��2&�f܊*h��wUah���䦛n��K����T�@�`~[p���nA�?'���eK5�6�Ч�yR֟r��.[�̲�8������;�\�J���>���;��|�n:�k�qD��"��w���՗�n��F] X�X�����$�)n{N�l"��tE0�6N �̘׿�m��RM�-��*�28�]
��#�$��|4�ew*]S=� R1��B�3��0��V��!H��ޅ�S=}͇w�x! �P�RtLi�c#���ޤ$���j�I'��4A���?'�4�� �P����:��q~��~}>�ʗu[��x����b�Y1�2|@r���2]tP����	���к�u�E�{� ����/|�ʨ�	H���ʕ��yxý�d�Y�h�����;.М�+����s,�����j�W_�Z=Ǌ+���v��V�m�3�fD�����ӧ����s2:��&bT*U=e�\q&fyX���� }+����I��,6Ӯ]�T@@; ��{��^��0�&:����l�@�|e�@�t&u��$Ԕk1��~���'^>�rԴQN�<&)7���ՃYb��`��s�"��? ���PqO�ӵH��"�Зz`�0���T �� i�C��F.�0�Ɉ��9�8K4ɉ����,�KNͺZ?��.i��F)d� �8X�\�{ҵ���<7����ۥd�&�O���x(rK�.�7���կ~5{Z`���Ν?~�ȥ��m��='�4�n��lA^�a@�c:�1}��}�=���/����W;�0,���k�Z Ӟ�������g�%cVq�3jv��	(9T�l�riDjUg�� �3�j-@*��ɬ��^��T쟋��O�S�����MDs��K����[9t}�"���BA�cHtu��m"�����h���͂^
�ﯦ�W��UV<� 5����%��DA�v����Dh��T�sBp�v�g�����^@���MnR[	�,��-n<�%�y��$��[�&�̶K�G�;��y߼w
�����a,��If�gc}���+�}�ϡн�oTW.��ڵk����C'�w�Ճs ����~��R��}NX��Kh�@JQu5�ᾃ5��R��c��S��i���5sa.1����TN�xs���������� �����G�)Mgh�0����oD���h��Hjm�ק/�M�1�8��h?��f��>7_ǄC���Hۍr�c5���5��w�g.�CuL����!��(����
����gS#��S�o���#_��Pg)�4�S��8rt�(�ã
+h�M�L-�W�g���p5�����M��mj��NQ����Z6+Ǧ�RC��kƽ�p��a�C�>�ǴK6k�����L���%��O��
=���NS����}M� ��e�ݧf���W�������og+I�si�	�2:6,3zg9!��1Z��JM� O{�N���4��]2:R��+��KfΆy��4�R)#]��NW4ҷ��Ȁ/RM��/���1�!��W�*2!R:i���X�h�UW�}�&�d�%�.�OM�����2���̛�)դ�������	c�"恳��+ձ��s"�240���,p� ��F-�� �vL����W��uB�-���5�SH`��J��[T�@� X.元fi�����r26<�n������QAd���t��y�Mx0Ƥ4VԂ!
u��y���� ����|���V��H �:�<���$�BbO	���^�����تZ���x+��o�E�������[������;]W�����E�:�(�\a�޿��䆛n��R�6��4Ȏ];=�������e��Ŏo8K��B�L�o�ҘS��&�/�X�ם�>��%�Ok��j>{B��BӞ����cOl��O<N�֟z����K��]n8!���M�O�����)�y�n9��T���7���>�nL2���ju��
>Z�數Mls�4��B0��dұ�b��N�F�r�i,��1~�؛׮�;7�_�j3��+��(4m�<���������x�1�Z��,��9�|V�n�T��L!�'��Ouų(J(�Jj�D�%��1�����J��r���u�:DQi�Ϟ>|*rxG �>�|��?u���آ��B7���;S�=�x)�������~�2k�B�(��E�9�,��v�ˮ�a9��ӥ��[�d[�<-�7=%��yiFmߠi�bM��0�P�q������Wʖ�7��%-ꁦ72:��9�[4K�=cr����J\,��^zI6m��4�L���ze���C�c �yx�[���e��D�����[<���F͛+����is�7	�-��)t�E널�H�<���x���b���{��k��KP� �Xq�1Y'ra�Z�g'�Tݴ �\r��C.���X4FS��f,�mړw`Uſ����ܠL��-tfKe|��������b
^
�hjd��<�%Ō=ya@!���lJC��'?����}�,=l�<�н���!w��S��d��T�Ȃ�K�R�ʪU���/W�cht@�{�Y����'�i���������=�������'+^�����A��'?���~�+SJer�x���կ�E��Љ�tG�|�4�p�򗿬���1����?�o8G3��

ݲn�:y�Wz�(���3����w�� ��K;w�=�/�n�VՔ���)�zqc��-�1�7`�1e��%U ���6�H�1��z���l�dr�,��F�v�m�]�WoF{�jm�"z[�YhX5�a�k�E���;����d���3&�̝׿��qj7>g2�7��͚��{�Bb�ƍHϟ��.9��u�םr�-�r
�f�UK�\�]
/���s�=�Y�0Y3���Ɇh�QOWs�"���_�d���85nH��{�1NS^�����i�ٴy�j�k�>F�S�1{�cZN#t��-��"w�u�8�%,x��(?\<G}��@�lذA#�H�1V1��%����u�a�d8Y63�L��E����X^1���%$������w&�3�Vא
M=�ˠV���/�Ɯ��%��,��ze�PU������vR)�j�=R^�=�ŷ���yki���K p�iphX7�:��(7]�t&j���U�}�L?��u�?2�Ps��B���ه�d��{�ys溭�-��~��Y}�<�Ѓ�e���e4&�~�z'4f��pEQ�~�Q���~���.�ixƔ�M�;5i�D��	#��������G����n�3w�6MX�t��x���#%�Q��M7��Y���?��?V�����r饗*x2���
�Bї�a����k��ry>�b�����#��p�t��h���6�{ob%��묍�'}�04l�!��2&��(/>����%ya��̎T�U�3�xr���'��3�>�<';�������0S��rJJ��t���������MU*v/�C�&Y�$f ����Q�����5�X �:R������D�R��P�|���hm��×鱳fg�.��pX[8N��s�	���Oʏ�cy��-*l�u�����R=	�06R��z�t}�Qg;M��x≲b�2͂A:&�VKI�1�ǞxLn��V7)��0Y���DÒx�k^����|��؝��я~����.�H���!@��Ru���j�2�L./�<��|��߈����,��b)����3d=�:X5"NۥޞY280"w��^M�����ל�)���$�	��������f����K*�U��x
�?��<�V���w� + Up�A��|Je:�#a��Y6�-�h��m.c���R�h� w��m��;��"�}�yp��0�];�� �p���9��p���(bo�xޝ�~��/�����V�i�3�s���B��]�9�����a�͘5S-X(���v3�]��eǎ��s�7��n�219�D�Ϣ�|`��|,X��H�p�$�7p=Y�f��C�=��(\��	��)bQD��!M�+��^�i�t̠���z6ױ`����Yݕ�\
n����K*'�3��҇�/�dj2�/�
|�.oqQw�s�V�*�=�1�uTS
5S*Pl��gZ-y����>�O~��'��Q�뭷j���ɟ�7����"o�;�Lxf�32tː
�U�V�+�T�`�=�͛6�s��
��JeU��+|a_s~�������QGZ�x�	>$F�ˣ����;�駟�A=)����Ro���(s{Y�?�����%D�V���3�tG�ԑ�j:b����ݡ��s���q4{:=��u*�����4+Q�^��, �U!��u�⎫��X�`�)�RZ���L{��)���x�P-B_��Zw\{a�{\CP$�V�����i�v2-��
�\��tF`3n�v�&.�)�դ[ (��<?�W,�u�r�9x1�����~��T�����;��P�
�7�7
���}H���'u�m�7!]����e�6 ;�v(N���(�5֨�)�u��Ti�R�
��ct���2�[��3|b�KVPE���.0,>�>�я*C�������MM?�zDqd�"��Ͷ��m�����	���)��5�`�&�mj����}��
��_�����>���e�M@���C1W��+��̰V����;0+2D
������(�m�ʒhU�ձ�x�,f����$i2&N�TiV��Q����;�
|�����a��YP������K����BRp�"	�Z�/x��ʑ���u���ǫZ���p�=�oV����2e���#�1�1'��X���7n� �,lD,@��p��#$�+H�0գ��(��[�����ׯ��E0��[�'�֩E�X~c� Ўc�k��{*J�4g���Ƨ��Z�lJV�-?��#d��B������g��WŦ��*�����ݽ*[�`tP|��`��[�S3�ռ���4{@TX�v�=5��A�'�GsX���D� �{��+��)�Uů皏B�.���f#�i���u��g�惻�o<%M�o~���S߱���ޠ��WH�[|�����ˊT����R��~���?92a�����7��.�`7��CVӷ���$Qx�+ΕE��-*�?RG�"��K��G,j͚5��!��$ԠS�:g�&���I'�$K�,��<�ξ]z�]���F�3�=n��A������(�!g����y����{$v����kt�ӕf�(���\�!�P�nӑ���h؉�9�s2���qI~�1d�5TZ)�̮`�O�'h��8���K�����e�Ų�[c��/S&���b��[^����Jf��9\���1�w��}}����x���'1��Jd��] M����?�~Z����&�?iER��4U� ��?��UK%�&�'R}� �糀�����8���?1q��j9��3�x��`m�r����JVp�E�s" ���~V <|��u?P�������O����_��3И��5�-�	9��g���.����C��lAl���0�B,\ &���R��o�y��q�Zf�� ������1ל|��˞�:$���#�v�
���h��&/���od�=���2�aЗ!�HZ�E� ��v�*כ�[�xOt�C�h-
4SɁ��"d��פ�<Y���q�����cQG��e���n�p�?;��x�y�6���.� S�����/L�s&�SS�i�������:9�c�o���8��͟�b !(f���\b}pS��	;aj7�ĭ#Y�x���,�i#��=�8k���� f<@�bQ'��*���@{�>�V��z������RKK��o�
١�B����z\�`��7x4�kLW�:�dĠT��ֱ��!�ݟ|�ɒ&c��;��,$4�k�'
��-Ȅr���wr�;����O� �j�������>�A��7�U2��2a��%5������.K� QK�o!�9�,*�ֱ{O�ERs��x#�_�f��e��߇l��g�}���ek�a܆i�w�駱�t�A�̔?x3  ��IDAT�^b��YٴL2
�yR�d�N:;��e��K�Rq�!2ie��t��h;tY�	�;����e��{A��B�;��ĽMal����g�F��_��EAPW�gQ�2�%��w��V|��hL{�?��'��(%w���b��	Q.U�HWf�T��er��q���S�b���Q۲B�fh�o��-)�*���2��)u�XF=�9��ŜC1�=dD��itD�*�cΧ5O	�^����5�r
!�J���w-ܝ�m����):^�Y��Vp6Ef�6��rkѻ$�Sѻ��lΤ��9�c�y�f���oM*(��1?2,e2)_���	+�5��;\3͘';e1œ~ ���uL���je|FQ��3
N��P-���F�* ����;����K����ɂ�L���+�?,]C��	���e�<V���A)� ��|�7�r|A*���3~�<�fn���$b~���Iiyu�7�@g��bE+q��2����hS�#�[m��G�Ķ����ٱ�������?������}t��� 
�f,)�fY�(�R��|j�A�B�C
̠�3kQF�z.�&��B���|�)�L��g�5{����m=L&?66o\\{FO�2�z���H�g��}���̦Y@6�+LE�ء�Z�z��`�z�S�����l�;d�螱��{�8��Ne��:���;�7v��9IE-3٨[w</P6�b���B9T�#V�/m[.M�ާ=�o��s���DE�:��A#�#��/>L����64]wf]��m?�mMlLl�v&�mۙ�v&�m��}�u��9g��]�]]���[g�֨ ���p�Z�+(i���Tߖȥ G�M�qdM��2�0'��^:x7-��R�af$eS�[���"*D_٢U����	�&uj9ad-Gv%N(BJ�J����
�ǎ��B�wh[��zZ'.u	3��c$��6:qd�l��&�%�#^��V�z��˚93�ٷ���g��Sq|ܥ	���ʦ�&�8Iz-/@<2��TG���<�߬[��X�j�jZ��U�������q~y�J4C��h��"]�j����R{rU�R��4ǣ����T��9��w�Ļ��<q�;�F^���.������LT�"� =����<4ƙ��+�����"�+1�>��T��$-�*��y�D5Vr�{�l�:�r�Ԋ±�Ey&�����1��d� u���b>�ѐ�N/�7AaU��R��o�tY1�7㻇X���pNcf�Ov>6��þ�p��wH�\��lI�`��I4�+�=�J��!p���s��ɰ�F��X8E�8�SԞ0o3Ĳ;(�w$�J�0�'�%v���
������ 9�:Lf�Wew���c)����p�"Ϟ�Ê����Xag�5&A�H�� !O=,��{�s�Лπ��.�ga#6�J�	���������-�%qH>Z���ϗ0_rP���R��٣�!��H�֛�P�E���7>�ic�����v��:w�:�I$W�kj�o�*w�[vq{��ͼDM(��ʗy(�S�}.�AO�?�p�����i2 X��MB`<���P9:�1o�}0h����6wp �4�\t]Q��@
&uUS:F��f�fD�*��y��Q�y�kSnq_�W$p�^�����Q��R����^�_�<q_�e�}�B	���N�o[3��!#b��V��.�e���	�Ȋ����~��e.�a$�j�\k�����l:�a�K�8���d�X��y��e���s���	$X��D����Y��S���p�?��B�i�)��F���Y�*
P`:RQh���e>��!�mN8�Ev��q��B6�~#����3�-F��������2�������ҟ� �R��U^��~�+�^?p�������濑B�����ݗ��o˂Y�Ws.a�J�b�Q�hT��'�]��M36�U��4C�'G���{wj��r��F���!`u����y��)U���>�a;����f#���UԚ�H6�뎛*S%�;ڼ<��3�Y<K�6��������C򬷟���d�=w͌�c����b��e��q�(_��1'@'>+�>�]�@���m2�ΜY���c*�x�z��T�S嘎���Me���Od��3ǔ���˭:h�l��1O�k%��S�:��쬧��SZ�ݾ�]?����S�ܽ�E�/�	�\4�M1��6_y���d�j���Ue1���ѐ��Z���,�j+b�4W��d�aɞ���D�����qAL\K��_@�q���s��Zn02��k�4�\�k��<6̵���[+&�$� �>���k�������� wf�:�V��>\�e���x�����*�;�M����F��g��K��;Lyk�����Fe+� 5iQ��.����4�������/1����Yj�4n*�����u*�֐��P�ɿ����w{�����ϒiF�7?=�h��.�bW:��Z��.�� ��U���ˬ1�x����Y���Ԣ
�W�ߤzB=Y�B�^_{��9|vڤ���%LuyU�e �-r��Jڷ���n����(�8��rk6��q�Aec�\�L���o�*��DP�m&O{y۹�o����8�3���Bi�H�~��P9�������/�*����3�%�#nR��ViӞ^0g�>D��,e�T�}�:�9�i,&y2��^�8x�d���4U�pQ�0��8a}�K��``������F[�2c�K�QW�n?���9�>�~?��nkw��-��������}_��}�8>�i���J�� +��L�=c
�+�X �kdw�4-�
ʘ��9I�b?F&�s��ל��本�">�IoL检�*Q�[|�ɖ����c����8�&,G��d�}wJ5
	;�#���q��t�� ��{�P��w�-a澜U�� ��@	���?z�˸KN�|�}���͜VK_�Q���?����ZE��~��}�6[���f�f��ߟ��U��0Wv���c��Ev��Q�	�YH�"�W&�W�B�xc�����RkV5�-��x���������z͊9[w�<����e�|Pi���R�<��q*�,p��*6�n������&��R��q�
�v�s�z�q��=�Uv��u��\�'�������i�H@7���I����ӱR�V�֋���q�$�+�Sw98H�t"�y���ݳ�|�@�ٴ�p�+Ŗ���P���u�m������Xzl���Jp�� ��B�m���=%����:��"������&k,4�}c��I KW���Y1�dx�O�ϓ��zM�>�zUn�Hv��/x�6�XE��S9�	O,�����PP"��i���(BZH�]l�n�"�Pnr0�i���b�o��$�Ѡ�j�Q���T��.��Ѵm�~�1>E��浱se�2^��$��w1��P�h2�Dt�oh6y��:ltL�3}P��<2����t�	�/��N�(��#x�bL�����Q��?0RI~U��?&[g�3A�� �M_F�I}7F���}a�A[m�/���ؠ�p��o�qD6-"'�_��t�_O�ze��sT�妅�t[ބ���؂v��~`��Pq�)�)��&�鄲�~�2-5ڐ�# ߫�D[��QH0�P��e~�Vy�I��C-�L��Lnk�6�a��s�7��}օX3o���b>UY�3}ف�u��ߟ�V� ްU{���@w���C�t��t^��w�*�gH���Y{iǑ0�\��~X��6�:��!�_6[�Օ3<'lߌ��>���'X�&Yy�4xOʕ�5�M�iDc���`���k�`�0qA	�7 ����I0@��w@@���'3��: �D��q6Ap��uX��R,�7qş� �N�����9{	#v$)�8���Z*��s� �������=�[�9�[yK/]���ZI����.D�܂K6�M3��,��r��G�X@lv]��.˹]f�S��T��,E�pQxོ͕K�m�'o�;7��\�1!2z_w�lN��������� ��&����v[�a����Ƀ��
�d��-J�����,�vUP�?�Av'���/-S0d�����l�2K�A�ړ���u�N�咕���N(����j]���O+"٧6�<�O�7��$ޝ���L���,^!=60��E�9��}���agM��%�O�4���b�ˁ�^b�H�{
P눻�#����v>iX3��#W�^3�_I��r���I�6�lc�����p��n�2��v�����4(i�n�d�N�ˢ�3ރ��+���Ӏ��řp.p���c3�]�b��]�5\'0���ۦ3�C.CS�k�[Ҋ(>{O�&1t�/��ȹ��f�{5'���Ϛ&h&���o�^[,.g�t4���?�cbm�P�%����X��'��ۧ�)z��
��7^��?�{�S?w�)LК�;Q:�3�z:,�13،J�toI�J���{7&1Y?���=�����%1�ޡ���V�p��Vè��M@����8��_����A�V�F)�ĸ�ު^�WՑ���*�.ܙ��h��c��|���DlJ�S}Π��ӊ����?m��,���T�&�%����������{�N�m���#_@Gc�ΙA%x�����6ɸ2���
�e�;���,��u�2庫���������~a�/x�IMyHvVb9�6�^��̨(\��O|�*���t'�l��U���=Y��?��P8g����^i?�o�Xy��3�"aZƟ;XGT-Z}����wy�f�o�侓-��Mq��lL0�R6d	�_�V��1$���i�c�OB�0a��� @b���2 ���i~*1���/�/I�M{�����O��_�y<?�xJ-DP�����qrb�G�ǂ�������:0��D6�:($�#���%X=�il	q��%���}U=�MG*/�~?�.�WQ���^w=��,��$*(?���.�����!Dq�*��NI�<��]�ǥ�T�8�7,F�i�����\�W��x^���+7{&����<�`��;@#��Ϯ�,h�/�s���K@��e���I�6U]E-�pj��a�58^$[-�3��.��e�$�������!ѫ�l�hO��91[=պ���\l�&@�u�2� %?�DX�s���bYow�����H��i��l�">V����B
�+0�[�GAKI8	�m�[�@�Q�̈́�X:Z�X#�O|B�@X�^���xwh��!M���E�q�QAsJo�e/гInv�{�������a�(Wi�5�>ig����}M:��=��b���W>�����Є�De����+TǇ�	t>;6�y��l9�F��v�6�������W$J^7K�W���`!r�Q}��%��ƶA�� �q[���� �A���M)�]�j�v���C�ڂ����ې�oS���bg7���C��|�خJ��}�h�=u?�.�E����Sr��T�ݸ*{�ݿ�%<:j�ܹ�o1i�y~5�Uq�d�D��kf���_�rAc�����śᅟT���I�}�a&|0e����?�6WN�t_Flr����1�y���?��(��f6�����7�[l�Gr#
��I+7� �Vk2~����L)��z�EG���x��W�Ӡ�~l ?�-ؕ(����Η����2"�2���ԩ��a�������(�Q�ffe�A1,�f��yj�a���5F�j=���^�ŃS�_����{|��ҎOj/ ���=�p�6�4ͫ�B�+ͬ�`��[q�MR�Z���S��gt}u�|X��2šT�W���#>� I�C�v�-�r��l'O��__q6V���N����Gw��1��x�����y���pP�Ӝ�鞐��ogiVģ�A`ZڻJ7�8��z^���H`�L74|������6E�P���GJ>DJ/\~6�]M|]`2P���q8T���lF}>�g�����6ZlFe��M�2�´�뿁�g��c�����Tڽ�z^�������s,�����|2��/
 >0�����mp��D��V���#4������ G��4�	�iC��Ԓ��tR�L������P�"�
S���ڷ�ڕ�&��<'�����{�c���t��ð.���Y2C��+r%̇�f�<�0/c����k����և���� E/-F&Pɫ�{:G�ifm�T]/����$_#��s�lBi�[��^���R�Eb$ZiF�(�#�TD�4x��F*�$�����p}��R��k�X���n��E�Gs�w҆�<���=��͚��;����e}Z���#̾�!4���)���	p<�v�0K&��\�M"G]Z���gf��?����%���7`h��.�P����m�ҵ�}v~���B�4�����Wg5���g��|6<�f_�=�i�;Ё�t`W8`}�� ����Y�۝���^f xsL�=��Y:��W�/�2햌nr�r�w���R�A�[���T�b6N�m�X>�6�.}|q�Εf��MPl�O�+�Y���R�oQ�l�U�.�H�����!8�'Fͼ"�EC����)@K֓��lY���q��H���;�^�r?+��/<տ	>Oěb ���i`�n @����`�!X�~�AFepB�04<7H���Fh�ܼ�iC���$�o��0*B`��oScU�<�K�*��8�B��Gi��'{�"��ί�+&B���V�`�j�����& Ͻi��*+�|���4e9��4a|�����������93D��;s�*-9Uܳ���$P�O�����*ίv���!��?V-:Dq�y�0�O�G�<@_>�nyo�X��D`;\L�9����xQۂ}�;T~��V@�(��4�ܰk�>��T)��1��?8kMi��Z8?A����y�D�!8�M푕�4����s�2��29�3L{>��q��3}z����8�-��L�Y=��@>�d�Eq=�BZA\\�s�;2�Zqbc�\�N�^ՃC�.�r�X��&\��ό��Q��@Eg�����DW���+!$1��P�O��9��ʟ���	����q7yi�u"���53Сz�����bs��U�:�sb,���˘\��W����!�{?5��c���Sc��y�:[>��4��Jg)�l��
�M�r���(�����&��b�@2�33�͠Q�Y���!��U����e/�\3@z[�5��4�+��MUnw/>��J�\IY�׃��z6E9<�F}ŭ���2K
��?
_��������#�lfE� #�k�^�7�&u�-�A�{5�{�ߞ�**��rI�$;=;�V�,��Z� F��/Pd@��<��6T����w��p� ���=���)�h�����'�3ٴNr�d��8=}�����Ue����?����k��t������G~�@�`;}a��){พ2ki.�R|[-,z�0�V���ex��/�2{��.D`�6��t�G�.��?ו����&$$�(2���M��l���O��2%<y~�,�s�I�i��;:d쫮C���[(�O9��KW����@�Ԛ�ݫy3nd\`��@�!V��>�XT~p�uá}sam���!*��F�� �B��2.���l��,��ȋ ��§[�7�~�YD���yj��Xn��Q��Z��ct
U׈��.�^S�g?/E����}%�	F��z������z�:���8�A7�Wg��2ݗ�E������d1z���T��(e4�#���\��a��쬧�<�~�Rٞ0e;6>�cO�8	����f ��:�y5X�R9��[ۜ?�%P�}�/�ҋ�	�Ve��]�t��!Xգ�[c�����k���!�th��c\m��	�EE�f��v��2G�R���5�1�π�vR
KJV�&2115K�T]Ϭ#I�������O��PRel1�&�On��N@c�ZcI�)���J�6��e���)��l��"�H�T�Q�V6�`ɼ&����A#��e6�!���<����Q�&;g��X��X�P*�+��˳"FOX�+��b�!L���Րd����(������p�G�.3�Uƌ�0T#f�/v�9�թ��0��|�����^+
���ud�]�,�)z�BOG���^��%y�=��'����i��u߅�*�:���1�i�ŝ�J�Tń����6 D���@�Y����&����+��(������� ����3�������L��DO�%+�½d�W�}R3;c�=2V�|��[���
�c�.�yf�B�BK-�X�А�s��s�+����MF��P����!NK�B������x�T�aӠ�Zbsݞ��:��e�%�;4�p_�v�0��ÍH�X�U���{�pa�jbi#_��	RԩybN����N�H�߼�y���"2��V���ui_�����k�X�]j8��w������F��~j{і����5��Ԅylze�S�{�P�P�9q��x�ۦ��Ɉ��ᶉ�ځhP����8\���j3g�K�c.G��h3�*W�a-W�&˦��/a-�Ȃqm~��CBZ��f�k�⦩E�5�A��10��h��&��!S��q|���t:5Lh�<8���P!�vxӻ��U]{�y�7����ЩyI��k+�&u��o�f݀��,���41�����;U����˴)9�q�1g���?��R��8a1C]����^?a�˶�� 6����WMDA؂�֟Ɲ�-�E"�W������������Ǿ�8�:��=���i�o���������|ʩ��'��,�vz�`s�(�J|lG)��џ�|u\�S��2����l������r���#.[�m9�<��%&(f���]�"#<R��o��X��1�ϥ8}�_'Mf�7��G�M�ƌ��j����*s�PR"3��	r��S��m���X����7��+���3SbV�	{ ��+
�fN��v���/�����/ΐ��Wl����SOP��_��|�)�ف���+t ��'m;�W����Ԕ'[Z���ο��h������)g�,Or�}}����~�]D?��+�fu�'���R������t���lን���< P��k"��i����jND�����$8oњ��ǐ��a��{r���r=�r�!��N���� ��Z��=�'�	��7À�x��vs&u,�Ѓ@��w����VʀS���N�)���V�h��d�C"�ĭ���m����y�7�@�N;��G����(�P�*Ćh�L��6�������;$����ʢ$�;�K�2g~�D�\�qUu�p|�*Q�]�5��8�	D����o�Yf?=gD_S�o�	΋ꮇؘ���O3&2Vi(��:+u$3��&�ځi������h���"vA'�}~,���sݏ�3�!��0����l���Eٌ����]&�9Xq�$f�]���h9`rM3�1��l6Ĉ� Pʔy����(PW[ n����u���m:6;f�q���7�0 ���B���F#�e_L#-����414.�sZ���0֙�`������VWd����kc��N�vӜ�x���
���z{Ðn�R�ya�qE%��r��q�}�,���L�j�"W<(�U��~�]�giդ4*�Wo<k�~��E+NР�g�>b�f,O������c� <�X���� į[�ѭ���1#~	ڞC��x&����{�M��	
&�d�|%�@'���^̞���"�!�|5 �	����V��y�z<�(kN�jj��p��>��`\ g�r��%�A ���y+nM�F���|.���{�I�L�-S�l�%z2a�d�f<��ǋ�<�QxY�	�%�'dn�K�-�P����֏j3�q�g�2ܿ��Y���1ط�Ƈ����#��ʻ���C:f�+ڶ�5+��C�H�ge��������}Vai���j�@ݤ�|Aw�q��K��Ҝ54&�ɣ�����)N5������{����4m�g��(`X�~r�H�H�\�����S��+P�4��ЉhM@��N�*&��o`��L�YB�����b���M5���"��׶�Ҝ��":�� u�'��[U`�_^��>_f�U���\�,V��������}Yu[
�g����a[?7��n������n�r#������F��ϣٮ[D-�O4�'j����9�^�E�O���:mwHeKB:�J�']#��e�	-yGK���I���yg�dm�9z�K'�x�����,<�t����1G�؆OE����2�:�Tj"99bDE�w������m�f��m˳���_m��1�1��Z���G<�@{kK�
.Ԩ�Eۼw�d�ctɾ��%pƃ�b�~Y�WTk��-c��
ED󰘆ou�2��]צ#*�QVK0����b-��*I1Ê	�r�+�i��1M�
9rU�hL8;�;٫�����c�^��ȴ��������a���(�}�FEiAE��h�3k�����faF���M7��Y����|�,B���)>�^�E�sU0�1_�	qrݴC�!�o��Z�2�%GRs]5/�X�]F�&>�����AX�M���g��P����[��:?3YLt���:vH{��R �C�b=%VQ��sa�^X�<U!��a�o�c������9��3��6w8v�"�Q(�\�B*�V6�\y:�ߗ�#M�o��4�>���ګ> �څf��� �����k��^����MW���p�N߸��n����A��Z#����8���ԨbFFn��mR�y�W�ǵGA� �}`���N�q�R*���L'5U,�ċW�L�ZiM��wծ#N�|���f��*�j8���ru���g�����ɚ��T>n�\��;u����q	��Ǆ[���_0FZm0��K���	���:EH�Y�G@�O����]=_���T���m�r2Z(zz�(E����>��ִ�o쨈�U�*���B ��[�lk��r4�-?��t��8�o��+'z�C_<�3�� ~@t����eveP��Ui؊#�;��B몀�^�-��Y7�:~<_G�E�*+�j4�G������s�~}r5�A� sq��z�������[��I�c�!�vhJ�����R�B�4��@G�c"�f.l�����jUbA��ݱM�����hz��ǧz�t�E��醧�N8p�!���ud��s4*�}"��b�Y<�6�S��`�����$C�(�JV�#�QD��e�TG=���W}P��tڼ�����&q���u��>�&��ڞ��dY+�|�)����&�D�_�4�L�Ԇ��9{��k��'D�	+ۼ��4����0�~��hd�u���g�{����xD�w���`j���0�(��~�޴y�Cˡ�ތ�#�w8B��!q�>X,ލ�Vz��������O�V�P���v����5�x�ٔo�rY ��&%d��X�qm/4#�PԤ[�����������K�~�V���a ��%��f��f�l�y���g��Σ��TR�gE�.�m��-�)���M�u�w��Ix�+�*��l�+�iSD>{=f�X�
/f���V����#���Ql�>���6��j0��5h��E�~��a�����z�W�����M�f{ݪ�JL�tqp+wK��]��觰�:m����2p�H1�q!s�3!9�����u�y�k�/��XZ,s_���|��Jʋ�k]5!�8�`�e�Ì����b:��~'��Nu����ʍ�ڻ�(D�
�8�x��܏�G����U��J�Fa	4j�i�`����1�L�f�P�Z�YOxĘ�B'�?���,��S�D2HR-�_���0�����a�F����jn;�r��~ʊ�Y?�Pފ��#�J�&����pe�� I8oo4MkRp�;�4��,��S���ͪ���l�����Ѭ\ ���Tc�H̦9+�R'շ7�����8���Ź��A����A�2(���F�\�;��!�4��ܯ�܋q�O�%VR�i&��!1D���~+��z�9���i���j9��_����V��0K�<�3[�9[����� L0���q�r(ڷ�m<t�φ5�=�!P��(gN�^*F����d�GN6ĺ演�Q����w˧�ޏ�j�Ӷ�Q���4�ph�L ��	��w��1����ݝ��"��.Y���$UL�R����O6߸@�=����X�˖F��@���R�!u��v�+� ��x2���(���g�͸ �qZ��P��8�	ru���-�#���~�#>��3�jC&2�@ӟGv�C��lV�w>����5UM,��+�4�M�`�h��R���4���..�I0f�?�,nT�ϖ�>4�[�<x?��}G�%U���0�D��0=馒����Y�4��t�lF������ ��k2R�Ԥ�^����GV�~���O�'�Ŗȁ{`������?=4�RzخAI����\ZCEj�ϔKϡ���_�sUX�$=�]�>;nfQoP���({��܀�l�H��՛�w���o�&��_�Aq�[�н�Iݟ��kxG����wi����F�B��KIh�o�S�Fo�����q�7xz[r�{k�˻N���@wN˂�+{q���Oui&��*ٸt#�LpŬ/���L�5���W��xبN;�W�n�'��*̗���֞�����1�*�ZnUt�h�ZӰ/ǳ
��/R� ������P$Ɋ���d�f��,K��Hj��Ll�rQp��:69������gi�c/̷�Z��K4*S�uוp	�땮qY�}kϛ���:���dD	l@g���#��E�fq��Tύq�s����KU'(���Q$��t�zws�"oh׉��F(V�MC��x��j����+Ȗ���5�j����?s����hu�,�0���=��\}=��d�
�c)>�&�����d�칤�]mҐxc^��V/tE��}t���aT�gn��~���kͪ��`����X����h��|��QGb�{9����E���cE�Z=�U�����Ø�C�C�e���K���k�0"6�d�}hʱ�}��5u��TǕ��G��\��A��K]��=��h�]�l�E�[_1+��Re�Z�ݢ�]ã�m=�]�,���
��]|l�coyiJl��	ǖ�1�VN+E����;�7$��٣#�&��`J�!bh�^���`�����IlW�0���W�3�ƺ/��q�b햢��ũ:<�MS�I��os���L����qFv��~���aDmlp:�Sۊ�pU�0���U���W�NC�d�t>I,�ě�����j��usi�O3a�1�j��gc�Z�Y�y�9c�U��mh�!�7 R�e��v��W*��<���滻J��\FrR���b/U�����*d]g��M�B(�K���L������s��'�(�A��&��=�����G��_ys���S��rW5�]+���e�J>��vI��.��MJ͒JM���F*R���[���f��+d,|Qee�B/��=kx�]���`Ѫ���9��uCX߅��k1���-y~�%k}�=�@�x�!p9�g��=��́���!��`�����'瓮�_�x^�o��@��'ұ;�u�D�oxS�rY�k�0%�g�^��>�h��=�#.U��_ay4�}��R��F?�J���}��rq�D3�BN�:���[��$���o�E�����&��d ���s�z.�7,"��������Ie�9��J2�fqLR��ņ�&�:�E��{���3ב�*���ĭJC/]��fd;��,J���\���
�5����{O�H�%>�O5���ҁA+�m�mB�8$�4�e�*}�j+�)����{��s����g�y���7��r=�z�S���pl�rϭy�z�#�׻F���[/�/f���R��m9[s-&�1��/R�%��l9�D���%
h��e۰#�u�kB��t�reM}[x5)q� '���sGӵo��R�n�|��"��)�{��;$Ӷq�m�c�Y_A���F������k��v���O�nxLg�m����"�3�*1�Z a:���I{�L��Y���kX�5���-�b	�	܃44�R�<R�׻�4؞�G_������#��͉�a�;̘���l4�ݩs$��kͮɾ�o\��� KR����v��3T8D�m꫏�Akc��TE�n�u�}�@Y?��}�� y��Z�4��c�)MG�ї:���=\�c��J��eV�� Q�	r�뢞��UʥOs��꿼���.Еo���z����t&���9/G!GJE���$�cfb�t㻗��b�(���Nɧ{�L�²��$ط2\{��	X���<�8��C��1 ����J Q�L7u�_�n�3 d���C���ݻ6�:��:���0����<�K�x9��7����w�jZTn��&�9踰a��0����ǋ�T1�����@|���8ːy�[M�Y����g:V8ݿ�f��F��[��r[�G���p��軨�y��˷����QP�ˆ���mu�3&Bf���o��d���0\A�΄V�@Ƨ�����Ӓ̋>Hg(h���Xg2�ix���}DO�4m�x%�̌H�����]-�?�Idր:NPTP�\����5�l��ѠC�YC�?:����~ޠ����u��y�y�8�$�;�+D�8����c�a�(I�h�c�;��r(Gcs@�ĵ]�+���%�`�'�>�#��4ٮ��G=��h�W��Ψ���~�~kW$	�q��x��.��� �m
Q;�V4}��,Ű�;��j�*�*��K�I�����������?�X<s��(�v����ʻ�sBA|���1��oY��}�'m۷2��f�V7�43��X�m������R��y�{�tbh>�CG/DvP�C�M#��O�at��dy�N<�ȋ� "}���L}�0�)f�� ),��0:��6C�Ҵ�N�!i����Q���d-�ؒ��x&~..]R-��/��e.����b�[�E&+�{;۾s?	I7���#P�ߡp��'�{��;�~,`x������6&Vpg�F�����\Ы|f��3W��؀��n�il��Aư��b� �j���f��k��92F��.v���ya�#I�g��m��_�*�����P�ߕ��a�^<�89"�A~*��J_��bf�Qҧ)[�i�V�+3*�z��*O���2�r��y��m�i�<,��%�྿7�Po�`�1(��O-S/�X��v{�M�]sC�zw5���Yt+7*Hb�㾤2�À�O~ZЃ����m�>%/�ZyZTw)k������K������j6��~�~>��b�@'��35��hGAB���ß�r�k� ����N�h_D�~m�g�"�$\��\�/�A�I=���\Da+���������Z�W��%�ʕ^:�I9����ȷ3eE��6�lRҹH�@16�L$�P��Gn�?�W���kh2A�^�g��$x^7!�&�������� B�LjA<��"R{^y�<��<N�U2�z�Ê����ɚ[���V�~:+��}|w�1���_ݻlߜ�XY�B�#A�,�1���'?�I4�S֝��3#���}�ヶ��k��ֹ�E! �T��?Th�'�/b�]�����R�*Vx��T��uXB0o~ ¦q�"5M�ɫ��os������%�(�Y����FU�����/��y�r��DѢ�J~ �t�{=�^��$�	��#�_�� ��E�ơ7����ҽ��#�EFn�ɸ	z:RU�oxx��X�?�06�oZ,4p��XY��~���	
�Ӈy9�%HkĄϑk�O���79� ������eK	��!Reo��a�'[l�]"��%��$�(�)A:�%����9qRl�{l^,��<r�-_v%�R3�J��2�╌'U�Oבb[�G���8�
���7+�fء68�ɅĠ#)�B��2L�6e�R��}�>Q��"�V��g1G�3I0f߶�qݱ�Cς�c�7VOS���ŬM����cy��Y����!B���ɀ�1�1�����v�����ro�Tۧ�����\�4�Ut���֣�g?��?�����\#�>�9� {���K?����s�A�����`�r��u��� h8U���)n�Y�N����R�]h�*��*�L�+�m}5���+�_��%��*u���E��9F���y��a����L.z�Yu|2fͮ�A��&D4�Z#�)�<"��䌦����'�&�A��xX����oӑ���I�FB���������5��|��0zw	t��7�N�m�{�仐Z0Z���h_����;��w��`�G��T8�O��������rZ����c"i!X�����Du~�he|�T��d�E�3\������eۏ�K⫻i�g_���ޅ|�c���mqY���Ѵ�>�*8�qX�ȠZ�f�|*Ԁ����O1��Э��O&��qᅬ!�^f8 �b���]����00�xՈz&S�HmXkU��~���w0>%qP�U8Q�.��[�*<ބN�v�Y0���xdg�����4��#L�kh��.�4����#^=Q��6�
9 ��o��L,�ߙ	k[ͳ�Z���l�CIK��]��=�zN�V3L��<# �6����/}!�(�QN�R�Gj�4ǟ��n@��w2��
�,cջM� �cRxB�ݫ�,R#)��W�m�����}bu��s��(V���?	r̴%�=�1�n�&6K�_��ˆ�=�6��Q� ��0�����%XĒ`0!W�b����[��G�Ə��=�5=&��
���pL��}��a/���!�b���H���/(�('�,d<��hϏ8�0�b�2�ڶ&dݧޛ�s@T�H+�$,t��2K��G�X�^EMcFv��d&2ۂ�eYM�8ZI7=In�D���7,�'\KXŐ��qa�6�^���V���.s�Z���t˜S}�����@��#�b ߖ���it?�ca�cp�_�D��"Q0�Ӏ�*�DE˴���qA g��@��a��Z��Jd`�d�X
����bP�W�4�����2�!H������c(��hS��+Z3q�U����� w@��n����\OY�LADٔ[��fQ �L�Q���OU�2->�ӅvvW����4�T�X�Ey�۵�F�  �Z�v��V^���Y{����Wsº�����
��xd~CP����_��o��%�y�J��E���s��t�Iv�'z͍���f7����,A,��/���Dd(�AA��Z߂~�<&�D�%5��<��|&a�����`��]۠�2޲�y�t~j<�9~��G�?��!�9�Aa����@(�L	�~���g��:7L�/�����u
<
R���
$x3���y��Vt22���KVy}j���-[��p�p�1�Ⱥ�{X��֮;2��<�kj�nU��=�=ϩ]�O�m`�f[�n�]#��Eg��������wXc*�����!������#E���	���z�B�&�C`-!gT<R1 ��5��>���;�$�9x�+^a�������L�=�8�ą�llv���\�M��#�o��j]�!2�r��R�����G�M��N�`3#��f��M���|��ށ怍MYo}�rJ(�E� �α��T3L8��K_�R�`�6�5���aY�z���\*[<o5ptʔ�n8,�V<�%���_�<��4��7�:�vf����>�-�3r� �+{��m��͙�O���3[�G�-�G��jj���P���d{hƼ�E�r�adF8�9�}���۷��-74y_���}�Z�t{_Z�u�Mo�2	��]`�Lf���X��h�Vv�5��cc��z��|�� Z���B�O1AM��!�������P��[�/n��-�#��=�	N�t��!�ʱXt�1���!!�b�ϳ��*��k-Oc�m@$��!$��eW �to���ޏv��ɺs��/��pZoI�4�lr|4}w�W����񬍏��/����DBXR��{3�\����,��莴Ӈ�w�Y}")��	� ���Ζ'��{��~�j�P'��C��/��,Yk|���kr���it$��);�3=�り��[�¿��7��u:N��{���`/������$O��g�����=��cNGcA���:�l��5���Kq��|��ڱ���Vڐ�)�zc��}��!��s
�}AG��-��`�}�L���y>b��#.�����0"�0B.������9��KC��]��{P��W�rn?�!��7�e�gX'S�j�6h͵����*�{+c�����~���dm*��]����G��~��Ie̜Y���=z\���G��O"�/��iC1�\��U�����{p�~Z�>zZ�s戮�?fc�۝�99Ѱ�;��W������^ ���[y�,S�L�{���66���$ͫ��t/ɣL
��(�t\#��N^��K�FQ��=���	.���l'	��K;(6����l�F�;�jW�ȚfRV�&�~����g0�>�\;㌳|--_���~�/�Z��[=�����z�pݢ���Kie������<+=��/�'�x��=i�֘�x��~���i�G���k��u{�K/�3�8�'��LJ0^%6q�#�8>�h��y��z �\&kQ��9F���0�s�(x/�|��f�tfs�����+�'E�8�<		љD�0d��#�,�ى���Dƙ���	2}�����"h.�c]����'�*g�9����SXO\O�qRP�!�JO��ݺ�lw$���k֬����:A�48ɡL�v�u_K�`�v��Q+�j�Z�CIy�%,�q�fV�U�
��u�s��DY!���R�>b~���M�/��j�aOm|����$�������Z��{vϝ��ӛ��W��5�`�,�+���6=����;�\�4�^�[�'ּ"�g�y��Y��v��e�n�d�c�����Aa��Z���i�sɲ۽{�v<7f�z�o��N;ͅ<�:mv�8)��đ�O�=c��G}����SP��^h��bzc��a(��"E6&�D�+:^��oi^��
�J(K��<���{��X4�!�ň��D4}�<���P�U����,&������,�邔�o��	�$^5���=��g���V�В�[�K�,K�g��O�ã�+	҉�,ڪ������d�����7����[*��wK�Sʼ�bm{�(��L#sK�Z#����#���_�`4�~ޒ����lI�'á���NL5l|l�x����/��b�y�a�=>əg���9`�����F=��Sltt��4��v;��c�ϱIP?bc��aU|a�	�vW���^���y�l�&y�{��]�轉r �o��o�k�q%��_~���D)�S�_����z�������S �K�ySB�	�L�
D^�ޏ�:#�^�}��)&��K�Y��)DhH�9����~
$G��5�ZP����5�,}��r����j(�e�A���-]���E�7�9� `hi��p�+4iY�4���\�w��6>9���@s�.���|{����o[���M�Y�E�N�sK'.�c�ȹ^}�7/c��/��7��G{ ]�|�z{����y1��Fmْ��s�6Wp?���SN����8RJ���;��x��"��^��zp	E��&�k����㫛6=n'��Q�  Iԝ?6e��
o��+��	�V� ��!������+^��g�@�cA��Dt��3ͭd��1��s��`},IA�����;���nd53g��&�R�c<� :�,���{#<����^S���XF� ��^��cnH���J�f�zbI���z����FV§�,ٵI�Z�ɾ2'Tp�����xF�M{?aɲ�~��oM�=̓�H��MP4��BL��t�������[�P\�Z����˿��EO)O��}��=��ԭ�uĞ���C���ڱǮ��kץgٲ�RSHG��/������?��O�|9�c�Gy��]s�=����L{K�]�¿Y��I��o��>�����b=�١���1�oƴq�&���O�p�|�^m^�
����GP\w�u�pp�	��A��c�wdg7�e���)��i�,Y�9FPJ����`+�+�N�U�Gʇ��U%�c^�6wL ����v�9��>�����=|c��{��v�c>�l���";e�J���,�Z���w��$�̂�N.�'y%����+��!��'��K���=�c�-s��R�J�����h�t\XK�����+�}��;�<��_�U���߁��xd�>�{�;����Xc�'Ň	�Ï�pX:��k}�<���#�<˕����ֻ��kiM4m��U��bMD�g�߳k�E/�{�RK��N�/��/fN�&βɫU��M��L<15Tw#�*���~�!*7��]�C?��ُ������U�)������o~�uW6�V|x	��M�yC�K(F�����G e�g�}U��0�!�!(F8�KxpN>ˉs����j� ��x&h15��"ry-}R|�+X�E]P��-���پ!�)}���\��,K�VYe`iV��<@\*W���=͖F��e{���k���L^t0��̋�5�I���l`pvڵM��Gg<%2�.��b�l��̅�#HX��G�I[X�R�j�����x.�:�H�7�CN�����d-M�-}O�^�ٞeH�B�]�¿ԍ��*����X�: ����g7�p'����崨�_ZN�C�)�Sw�Kբ��Ұ�y�L=�gV��63������{��`�j�� ��m���C�6�K6Y���ñ��?��O��uϐU-Z]�dp�^�7��ω�zXj��y�!�����*՟s�z,�qy��g	l��ܛ�N�.���k�\�"8�S2��jȒ�a�wZ}����R^A���t:o١���cɫ~����d�[�:hO<��Tyi�HR,��Z�]���\�YO$܋�U��F�9w{�x���퓶eێ,�ײd��h�;7Hs)��%�!N<�g�<���c����ەQ���	JY���+�{/�rqT�Ȓe��z��}�6[�r�mٱ����X��?MvO�<�Mأ�<��Q�O�Y}hZ��41#Vo���I�Q�vȊ[�{ܶl��欳�*�Rzy*�Y,,=6���h�(h�U��%�����C�YA�K/����R�S~A�?C�y��emɲV�%����0�����<G)��ȸ��T4N�:k
1���m�g!l����E0Od�Ha�}����׾6S@�v{S���ط��9$3U���-��cTbw����{�/�R��ozf��6����$,���t/O��q��$�К�q����K�+��4�7���j'�u*���i%H�^�mS3�k_��~����!��!�0(š����S	���^����d��x\�5�j������������gmbr�ο�,[vH2PmԞ���m����M�:)�4�?����W�>�,b��|�N8~��%����`��w�m~v�'bd1�J	����$�e�~�!�iXlR�{UeѼ���׼�5E/-"ea�qם�����w�/���b���nk�^�\�1cFA�Nn~dIȃY�A�J��>:���]*��f�!Ų!�.�Z�*8'�qxZS|E �q~��
���.���u��攋��4#�gF�TBV�ٰFS �j*F�ߔ���>�{d���`�Y�9��\��_~V�� u�/��H��V 1�+��d�`(�����v�/���7���������=H&�u�]^:f�-v���m�s������� O�֬]jûFl鲕����;�زQ{�)'y�J�����{�"ٞ�w�V�|`
���/�������ڹ��V�X�A��?�v�x��ȳ��5�竖���O{�����t����n!)���f�����G�f�����ۋE<:8vHX��M�9<2���Z�I��Z����I�߼�< ,��2�ʊ%H1��t}X���Y7���i���~,�s�<M���m
�CP�9�
�P6 K���R!���� �(2V�q��hgҔ؞`��d�QnA0L��GP6��J���������B��[@!R:3ɽr� �m\ż�H���Y��{��
 ���y��fB��Տ��Gp�q��e�t�HoH�߿�6=�ɦ&F��Y5�Om�dK�bkWeW\v^:~m�%{��-�u�D��c��V���0�)�΃�~�;��;���68�o�#%;��b��m�=�̟&�1�S;����/��ի�M07�ζ�~���{��%�\�A ��x�^np�7���H��3�����CPV0�1�X*���rW�f;�uZ���`I#�# �sqNA>���'��Pք���
^T^�M�`
�F�c|�-�׃����HB�\^zd�]�Cu��$�"b4��HT5U��,����e��T:�j�2ku�Y�	b��
���\��_��@��h͕ 17����+#����}
멼6�!�Q̳�#5d�w��;~�*k��ǜh��%v����Ș=��öb�!�b�Jמ�^t�u�zOv���w�{]R��ҵ``�|X��?���ߦ�\���j؏�3_�o|��m�в���^}�v�k^�Y�XC�w+gk�0, ������X�:��l@(�#��f0-66�~i�}pt�hl`6�\|��W�R�� ���H��Њx�b%|q.� C���C�V�`����Q�]���cbd��^QQ1B���׃�y{H1Q�2��}��z�R�S
��5������x��&-�
�ߖ��
�>]h7m�׳�Sn��f��?�{�
Q��r� �4�����9�������x�}~��󁒅�)
hdW)��*����y���=j+Vn������7$I']���G���F���/����v�=^�F��}�.~��*���MF�ʕ�=SʉA�����ܶ���.��O~I�*��<0�ԅ���pM�5��޻��	"�N�j2�l(�?�я��� Y���{.��U�����V7�F��o}�L��_�Ln�R0@��ɳֹ�{�O��;b���� ,tq��W�0G(`�5BT� %֮����`ۇ�r�b&�cP\��(^��W�ҹ�%%a�V?�60���<R�5@���D����Kmf0�C@y=�v\K���;�tx)�������f}�|�H�-r �=���Tn�09<(]�9�F~^$L);/�9^��o;���]l�Y�k�C������u#6�d��عծ��Z��G7gl�ь-V��3�X�¿�h:elddgf���&�s��o?��v{��G�\
�أ�v�N�e$�fvo��6{���{,�F�SD�����?�C��h������KH0x������_��p�YXjxp,�P�U��SO=5#t����'�E#�폘?CBRyZ��Ǆ)�}h�cP] �t>����G���,�I�F�JHIgA������>Q,JTV��;:��l�{�<���e ;���ؙ?�Y��Z���]�ᡒ��l��{��b|y�f?.|N�X�>�6bM$����I�p>���"���gV�����x��<w��7��	���o�=���u��?~��vc�ݲ�5��!�n����o۾��ȕ(��G���4�����7�X�¿U�N�ECg���W+W������2͎����h��@ڠ�b�U�z@ic0�X]*��q��;������)AE`"(������2 8�`a������M&�Q���+P+H�y��3��$P	�ך`�F0 x���q|��W0v�S+�22��Jb�7V������J̍TO�Ž3��4�P�PD=�{�k��_�F���t�l<��P*,��&� �C� g��A��R#h9{�����,���m�pD~�1��1xy��{���+	�������A����	ni�3��k_��?+�Eo՘nb��ݶcǮ�HH߅g�{x��T�̳Ƣ��GZ�Su���H��#ɵ���0=�:����i4������d�Q.��=���ܥF��D��44�����C��O��Ii0�0��#���M��N�'V��KL@��|�`�`�tB[X�k�軕���=�ǜ	A&*��?����x\k�vQ/���:��(�I�3ޟ(��B&+�*�C,��;dH �r�:����J9w
�%�Z>
�b����l���P�]�>?��`l���<���i6
%��(XS�\�6��9y/���l�|9+�9W2W��Ox6q9�}��H�s�4ʘ+Z"��K1���z`�(N
7�����=�����q��栘�A���G����"T��0XC��Qʆ�c+}e9S=�S��J��l�����d�Q|�+��E���z��ڸ����"b��lŅ"�7�\��K�D���E����BK�Pcq2Q�|sV�s:�>�wxE
^
�%h�������l��#��m(kz	d+�h���E�b09���e�k>�<�%)��ȥ㣱 ����ܷ�T�,�u�NA���	���me4�y_��tEPˍ�z1z���3V#.�>/�@7�̸�*<s*�:-�ޚv]{;b�yUڧĀ����@�����1��`��=�{�̣R����{��E/�{|go=���:Ӛ��6��?�y���aU��� �������>p�c[m4-�H-�9��mp�Z��d��ǾЖ�(��k�z�k#d�=�Ȣ�A���	�U�G-9x�U�E�by���Cשu��v�ɳ�x�X-�	%Pe���B��!ڦbU�������*��"�\D�z2��s9�`�}�&���aȋ�E�m�Iq�kjgHO�=���sYM����ڰg)�c�՜^uS�o��ٵ�bn�*Y���y���g3��s���]3g�*F�gV���_��{4g��sE�\Q��C@������r6�,G~�{�.J^l�.�@�p�v��mp>��N(`(��B`b�r���c"�Y�);ݫ��7�����b��u������0�O|�^�G���m.���:�_��`4����r�3zF������3|�*��8A8�Y�4AN�֕
�EA$�&!��w�N~9,�}ҋ�O<+hܫ��")
	J�U�b�n�2%1��IyZ���htXx����{�}�D͌*]��_aD�b��wQ?�)�U`����^������(�p�	�qi�,��YQ��ͭ@��T6%���*�Å`.�bC��Ҩ'X����õ��׮T�,��χ�/Z�P���8��hY*Q}%��g(�B0	�/���S���΋*M�0�CL��9kPP�2�uY������Py�����0�C�`�x�:��T`�)I{gEC��P�Vre�r$�cs)<�K���>JvblԿ��#��ƾ�[�x��5��PW�\�}�'�۾랻3je���3��"�.���yD�;����l��!o�y���G/�f�8��6�bD���m�շSC�J�Q�`�K	6Zp��TS�H6�m����h������X��}uǠ����Z����9����{#���|
�	�ݟ�{�C�A@$zqR"�^),	�s�~�o5fU�k@h��#HBВbGz�N��ۇ���w_	y1�$�4���nCumtm�l��~V�.�1R#���l�[]���%̹�Q���L+y�*q+�F2���^�c����X�¿���L?�g�5�.�Y��̔�� WPM�{��e9�/�_~Yb����f=��n�%��X�,/p�a�~-��u���L��r�|׎�UU�.s��9O�%Bϟ �,8��g�u�c�	�^��ye5*CT8�����$o	+��V6��:�X&b�ț��8ߍU�^��"�7]�O�S�A��P�N���X�VJ���,"�:���n�R�i/��k428�k5g�Y�	���3�� �C����V��a|1�C���ǿ�س��L	�1��o�/{�m[3=���L��5���Fĕf�`�j�ֺ,5Yڰlq�%P}��zo�XbX�.��r�^
v�M�0�F�L���k�cD�������� Ās'�R����}|��T�-*{�C�,oi#{GX3��n��_�ñ�,)�5)%� Vf0�ٯ��
Q��x��̫n�W�)�:8/�'�*,~h��>�=�r�6���a���O#�Ә��i�hOkϪ+\�w]�n�gX��sؓs�\ا��nf��T(ɐM�H�|�g`��|�X��h�S��j�K�F�/��P.qt�5�����V[xE����,#]�R� ��\ӔM��H@ĎO�4v��=]C'��=Yt�0�|C|�j�p����eD;��g��֊���1�1� n�Ź8V5���9��5[��,~,v?�FLYE ��T�?*w5v���X�3i���"���nR�P �:c�X������in����U��e�4��_�1�O�gQ.�Oĩ��L��֥�2
}]���u龳}���~n�Cy>�d���6�!��"_ �����@E�^���}(�P�fV�X����f�)�x�q'dV�Ĥ�G�mٚg�V����%�!+�����Z�F
c''��-vX�q�j�+`k�hQw~N���3a�^�NX�ҧ�PbP�G���GB!2g����PB�y��+K�90����a%_͵ܶ�έ��3W醨�Y#@�
��<�	U�Gx2��O��ד>��se�F>�=q�W\qEf�4��`�S������z) )�+�9w�~�扌d 73A��׭�ViZޅ�����K���~R�=8_�z���'��1���^�-҃Y'�p�y��g��@V�i��K�����
`��V�'C�4��7N5	��1�:'/y�K���3���)�:�&��d�y���'K^�	.&.��O>�j��~{��fcSD
!�[����`Y1�Ŭͤ���)dU����GL#Y��F���QK�G&	#*3)C	����!O#&��߅V 
�I�<"�F�Ne�
��^P"�G�\
E]��1>7�^BZ��V�̺&���:G������JT��!��2�״6���:�����9���z
ȫ%�Kq�n�[�Qݓ�Kk�כ-���u�s��j�+�"3$�5�2���G��^��N8�=ϥK�����n_?��Ńv������lyY�9�t>p3|���U�gVOQOG����|�7\��H�HL��f��V��&k��u�i��op��L:�~��~�7��_���\i\{���]Dlu&�Lc�4{�N7d�kX��%������Ɋ��YC����Z�Ŏ����N��ڬ�.��(����u-<�d������,AS���z��u%���6��/(2zCR���o��0^BK]���u�μ�V�iD���T�UDl����Dh'Z�b��we�f���lC��O����~ �uZ��W��(���!&���d`R���3�p�oȕv53��9�l����䦧�_�G7 �U"�P	t_Ǣ�y	�YI!�Ed�j|/��"��񤝫e\�qۼ#�j�e98X�ɴAN9�$[�f�O�����ª�P��K�����|�7ۿ��������^�Sة�	Pa�sI�P	C_MA�� ���1K! ^��C�G�j)���'�
�ٯ�r�3v��,x���_��(���Θ��/
�s�]�ys�L��zI ꘨e`Ȼ�=d#D�s�L*Qu�����y]�	����n/?�ZPRН���Q�1`�ƺ֩F����Y�KAc=��&
\x5Z����4��a��⾋Ɣ<���Ø@���կ����J¨lN��(�8͂$���ڵӖ,�����>�[�/|�Kɀ�ϖ-Yj��#��q_Ǣ������˽�����^��+��9�H���n���Y�W�\�=8O?�,��<X)Z+^�	D)<��#>���_����|�#^��f,���� ?�5��׆CyQ%/C�v(�'�9��~�(9~t/j΢���5����lV,,e��������Q�Œ��$ "�����qi.��z�h�Ȑ0��=�/Z�<�JR�1�'��R*�������R��bs�H�t��Z�E%�EZ�s��'[U+E�YJ^�+���q�6"�罠���@m�7%�̟����c�~�^ӱm<\0��z��ב��нy	���0������R���7�>	~��~��6nz�n�����;}n���=�<[��P'�,Y:h�~���_����^��A��v[�¿Ճ�59Q�`��]#v�1G����d}�U�?�arٶ�q��Yv
��/�ݞ|�q;�e�Y��RW_|�G5jg!bI���p!I����ۇ?�a{����3ZGmj�|�6��(l�}"@X�����k\�h�	o]�g��9Z�q=>��X�jT@�8�\	&Q��[B^TG0N~7z�Xx��6*�X/E����xu�*1���u�־p`�S�]T�A�-���y=Blj���C�3&�˜0W�a���=�X�ū 2ǣ�E!U��FC�q�Z�_/��@�+��(
���e�����'wq-Y���;�1��3'W"(��<m۶=�s�C�����h��=�y�k�A%��g��w���2I {n�3v˭?���m鐕�%{��_�5�����^w���V��UW������vNI��Ƣ����dc��\ȍ��N��m|�Qk�ǒ��O�t�UrL��o�޴�׶l��w��}�ݑ D�M(�#��F�W4<�dY�
|F7�׈L�N�!��M��T�b�Y���М�sa��@8F��x��
�,S�	�X$���*!#Ꟛ���D�I�="^�Z�RFX��	<:���l7�' K[ޒ���.��_�3w�F���������q��3��U0a���jq]��՝{���7�!�-4�5�>��Ϻ��� �8���q��<��Ig������ܙ�+�?�
�zQE�������o�o�q���\��1��?�>�[�y=��Rԭ�1{v�S�s�6[���zkmbr��Z��}�����ˮx��AA�u�v��?rJ�/�K�3&��Y�kIz��^nL$��u߽ގ>v��o8̞����L�?ɽ��)�oO�J��Э?�Ņ��ظ��8{j㦢 ����)�.���B�_����n�tz	8Q��^GFE�5�G�g)XJ��\��,>5���*����BB%$T�����e&�@4Eᘂn�#��`�ApR�k��vX��/4癝3ǡ����i�iw&�u+w���Y�\�փ:o���v*�^�J=(ʔ�����&R�������|�yWp;��el(�4>9QԧaD�c�F��@�ր��+Z���״�bn���]�J��v:xql�O!�F�<CFRr����oذ�~�#u���o*�;��Uo}�-Zb_��W=��o
k�b�z�+���+�mz�qk��؉돰'7>��~��F&_���-�����V;�S�_���Jo��hvx��@�������;��;�V�\�&��I_���u�G���6�`�)X�� [��1�,(K���kXO?���@*��𖷼�q>�,����?m?���E@/�ᴐz�N�Yt�8{W���B� ��,�����o˞��>�@R���^�Ғ��+!
S�uH�I���|�>�];-���k�gAO,�p�^Z�zL�L�Z�+��|�[���gd�Ǻ2���	B�������&6̹+�r�5��	2�ٹƤf*lV.5�&�������A��KVt	k_�����s�X�b)
����?���Z+���~��N㦮����<�����{ϝ��C�@J@�S@E�����T� ƭ�2h��� qd�	':DM< ��g6�A��+Ib��v�����R�d�?��S��-�m�&3�Y�T�R���L��h7�@X
Fbc��	�b�}�;�q� |�w�w��?�)��Ul ыJ7pd��������H�0J���	�$�)��<�J����ıD#J���P��I��@4��D.��1"�U�
���+���������;Q���>fbGVH�̙�ye�:� �ǅ�G9K�k��(
�v>g����g�W+X'*9-�W���fce־_���ݳ�{+�L�]O��:��ÿć~x��n��!��e�ā~YGxyt��|k�����m���y�!i�ҟ���N��O�s��=���o��VK�x]�\Ǣ��L_���0D��rˊ��Ov�����I�*-��!��X�C8��t�y�{�:��ƥ�'-ߨ�N]{�L��@Y�)��ׁ���
03x��4���V=�$P�(�)I	+}w��kr���B�\��b�;RW�rHiʒ�	Uz��+��>���6��ˡ5֔<��{���k� �
d���?� /�Y�����%����,�)gP� a�
���Q.�z9Nީ�J�=�L[6� �`���c��BI,��3�bє�u�O>n�F,@�%�� �D���-PE��O�S��4��i}Y����<:�ÿ������OL+s�)�ۈ����i�>����l��z�ȏ9f��t#�+K"�L���db}9������H�Q�H���l �"�;�3N����Z�!��|���ǚ�lv�HmhY�F��1�����Y��7R�$@�����R�n�SѱN��G^�8�ԘG!J�1����������6S�������P�q�ְU���yMA^�Q�C8��"��d2�R�z�/(���oֺ�ː�I�����?��X�)L)��-TF�c���$���O�q���-�׫^~�S�K��p��ۿ�A�w���M��w�y������>�o�!���[Cs��_s!�m՛S6���Z��rr �ג���2���Ĩ�5�!f��9�E/�ͺ�wgg3`~�a�j�a�;�OѶZ�VV����Ln��'m�ݾ!�p�$&M�*�t~YbJ�<� �"ZR���lC�����`���q 1��6	l,D-N����q�����=���c�^��V]A��y��"�^����%mJ1pH���+Ȅ��f������^�g.�_�M=7��
ݕ��uQ2���Aq��0ψ��=A2~e�j]�X��o8Ya{�F#�k����xĠ�����i�=͵�Ѿ�Rkv�L���mHc��{�s���W�ʧ���8X~�m���<;�XO��������X�3C�������,����lt��ɦ�|��>gcim�Tdh�
�&E2�\�¿٣����l���^y�����s^�lOۮ��l�����F�(��Z�R[����a[w�R��#I�[�8�2�#�KO,�E1(
�ن,���`U�W�_�;���}T���X���r��bPL�t�$KV�
���A��C�Kx�*����v�������n�M*�D�LP������υ�h��f=��1��
��2�A�1j )���`p>QL���QS�L�Ab�b���s����]��cnj��r�v�ry�z��0�-�=�N�n1�00�{���!}�!;�%��3���۞�F�φ��:��4�v�I�أ�lLϻ�pF_2F�3��w�O�&����;��9�i��g.8��$�WZ�@5�W#���:�t�?�g�Ɇsp)�v��.*0m&���l0�?��?م^XP�b���G{���ͯ`�\��%p�0�YE���>��f�9����H��s(���C�0F֢��V\��͓!�\�AyX/�>�5<��"��h���6?���$%X��P�e�� �,ƙ���A����H!w
"�Oтǻ�F��Z;����C���ľ�,��̚��o��33��o�s��&�^�9��3��潔@l���-oՍ��z�a)~�'��7���>��[�;e0�&Ӽ�\u��ܽ+}~�m����J�犲�f�d�Ye�^v�{�z�<{�F�����/�Z����'�BIf�;��~�n��&��5�Nx��:f�/͝���'7�3<n�rՎ8�(;��uv�y'���MǺb�p��^z�M7��"�gS1�K��B8W���Eb)0���lB9&����|�7C��K��{D����uQ�-o"R�Ua�XH1��x��l�wO O-��cEHE�L	��6��Y�M���3R��m	r��P�;��g�a�8����D&�����W1�"~��dp>�����`�2�*�9���i���b^�_s=)�Z����z^ܭ4͢oN���\���zT��*ʹ���
쿈�NRӿ�����\�h�����/
�ꫯ����ﴖ�<;��+��,	�I[��4۹}�y�i72��ɲ">s\20/����~�	�������n�G~�ȍ�t�N���*�¿�G�Y0Z��ot,���K�y�?�X{��׻u����/�ڵ�rNu�l�L�S����X�r�� ���o���_��c�4��;X߸���o��"�3\�cb�	A+,D0bY��,�IٿwW����/���<#a؂��6�%Z$�*�~�И����?
��Y�<�'��7T3ch�ƫ��x��3mB�<X���_u��.R�,e�
�g�x�j��8֥�-1+���3��^�?�x�.�����Ox�bŚFsabE���B��B�%��J���L�dk[sR}�ݾG�K��BŖF+�q�Y){���m���Sݽ�^^����~eE�&`�}�_�ߏS�eyƬk%H*7C�c�Ĺ�/�ܾ��>�ev�y/�����)o��x����������lȊ�ױ�/�>�wı��Ѧ��g>�Y����� �v�����8*���6:Fᬺm߾���o�օ��ZL�����x���������.� ѧ>�)_���]��ψPL��Ŧ������ fHH��8� A�(PX��s��糲U�AHΏb�R���
���:�%���M���D�,T�AX�|��2�D%�
�1)�z��_��_�k/%ſ*PƘ�k-v��Ǫu�kS��
�	$�.a�3D)�9X�Ϫ�C�T�����JaP���_��`!�i��>A�F�!���"��`��H��9�%T�NtL�@5��`�:�t�&.������d��Y�ֱ��ã��̳ٺ�r���2�;STޑ�zŹx�=O����\��x�rX �7q�o��^%��K.��Q�s�)g�`�LN��̵>�����{F��j�k��V��_Gg@�QY����W�CP_p�Ey�⩂~���?�1woQ�E4K9Y0X����Q�෾�-�.��B/�@�@��
D�E��3,y0,BY�
؉��*E	E�D�Q�/����|��F��.=��r�=�C�"����@
�r��'b�,4��7j̑� L@����ΪT�EtI��Z�ipN�s�)���2�J��9�[��*!+[qU�d�c+P��c��cL`�!E�ʶܻ����c���x/�"&҈�(�]p~��'ltx�=���6�kGz�n�[��R�"@#W�<�,�Q돷#�8�cqO'��^zzs�-͗,�93�=�,�'��X����Po��@�-�l1��s�v�w��x��_�m���a�g񙆓���k�X��sN��?�Yͥ��q��/u���d��M�\饎�e�Ъm|j�mݶݾ���x���k4�%0>�Sݙ�����
�J(�E#�x��21�*( b��JP0*-�6�'˓E�LD%)H(]TQ����'�������#��Y"A�� )$��n���V(�eM�_�X�!���w�k�Ϝ��{|���3a�#`e�G�q���C�Q"�N����wz%��x��ށ��4Шp����5�Dzyg�\u}�A�ɱQ+7�WI�F_��+�Y�MU�-�D���X�]J
#c�4�mE��h�s)�/+�s~��l��r�AG�^�L���y��
2�JwH���o�F�G���xR����p���y*s��N�j#���x����e��RT�^�+YU$`d�{˃+�mg�wʭd�!�x��;�g�UC�e�C�^u�U�(O;�4�H���T���&�5r���| )��X�vK�ɢs#���d��'���|*=��Q�?�ѹ7�AX��? �]V��V�zY��k�J�Z�~��`���)� L^������)oa��TyS��UDN�[q<[�?XW*/�h�9��b�sC(���'��@&�kdl���wHA�
*l���E���~4�C�.���%i�٤��[�}W�fΓ���̠R��M���ʜ���{ �v����6��=���J@g>�|�W�*&�{docpѷ� �bzzf�ڱ?y��2�3Y�6=�%�S�!����݋�S{h�sT���g.̸R�t`Z��m�ˈuWD�t�%�_�k�� ���`���`�F<�k`�I������E���'?�Iߔ�A�p��?~-W,�����W�v&�)���,PY���c��|4�N� ת�c���`�^\R�����p�E�YpLE�8�0Q#m�K s�Yo�f��|.�iމw���L#�de%�u��iK��ol�+v�0�N\~=o�yQ�D�7oRק����T�X��x����p�u�0o��$�T�GU,X�s�%�e��X7F��l ��{s[�)7�j�	�d�I�yyh��@溪bB�AmdD�����y}��_�}N�7���������̟�nȐf��J_�&��V�Oϴ�ɣ��~�ûlp(y����ʔ 6��F�$���&K���6Z�"�~�E���f��d��m�z���K�1���R&,����� e! (���O���-n�IH�d��h�h}Ja��#��%oɲT0W�Q�'z�+�:f�"�x�AB���E� �K����0R�N�
��F0�@�R�Q)1
Aל�ZKi)�b&���<������H�a0�7��%�5=	 ֔�y�����l#�1⻕�a�r���I!���g#�-r���X\�ۂ�Ӝ�f�Y�i�%%�%~a�;%t2p}U��t~�Ԫ��!*�8�W^��ɑ<!ŋX׼Ϗg�潒�HX@`��dՍ��'m`{��J�V�Z���I(Zg2L���Қ�� ��}5�x���du��Cm�ܵ,{i��H��Rő4��0�O����[9_p�^��w�>������M�{d�S�c�,�����˳keMŠ��T HG�B��x��rs�Yd[%�D�dh�r܇(�x*׀`'\�d�q�QF��D��7�hΫz4�.bYDG*cy��[FgPS��C}�f�u3�ۿ��΍����s����<+�*q� ����ׯ/�S�]�j��bs
&� �G��<)��R"XΚq6K~OJ��[�E\ks�,b,"Χ��2�ߨ߇ ���N�C�VL��<MQm�3�۩�1���<��|��6F��~��Y�H}���+�$x�PQ��<��QfK���0�־A��\��G^�d��3{�g���y������_,�i*��^|��2�a����^_0L',"�}ڵ�r������z,��c�,LYw�?`���>���x�*� �BP����[��#�&��,J���Hu�`�}�m�y�G�x�l��1"J�P̭�%�n���@���8V����͛zK��,TxO��I�L��Qָ�4t����Cl.�A�~���$�8�g*�=�f#)����ߏP�{E�¸)&#o&��ϕ���܇��R�ϲ���D�p~]��}���o~ӫ���?�q��C?���eĐ��׬C�劯!�F�}��1z����ح�0�j@��EL9��큪�k���/��/�ܲC��h���;d9��Դ���zt�&�F<9v������mL�(j�oh��Q�H���΋�#.f�
��&P�Y׫�$�#g_�X�F�'���{���s&�G���*X-���P�^��+Y[H��!K�&^��Y�xK(�X�ZZ��-?x(O�q*)A^S�G,I0SPV����-Ԑ��<f�S4�͖�"���ͽ���*�`����-'k�Y�y��5���%zp{��kDa��%(��vT�Z�>�`1����6<�*��Zӕ���j�i,k��f2�H���HY��}/�r`F��e){������Y<\�@PDw�!�u^4%ܦg��R�����9GW<ZȲ��Q��b���$���~���K(�]�ML:k��_���;��$�:�[c�}_�sӼ�p��7�SA���@y�E���yw>/A"��WF�^cJTQi���s�j:�֞����4�߹���ӳ�wLcy%�G�n=�z#=���*"��6K�P�-*W�,�w�`�����<:��)���Bs~���x��PL��D�P��zS��s�[ƙ���dzɍ�"�n�1�:iN��|��¿���5���6y�	(հ�ZY<�'�]�/��z����fV�g�D	�J�m1���[�i"�:V,�SP�S��'���}ˊτW5�κ?1o�㗒yH�JTN��,��Y�m����ڟ�=�OV���b���)�d1���O|��1�S<��D�%�y���He��;��G'$ة����^�������b�u�T��'w`b�&Y��$k�{�f]�X_{&y1��z#�1�ǲ� � ��ڂ�<�k��;h>y�R��baC`��@�xn������9�Cc/0�����F/2����,��=���X�¿�m�6��$,�k?:U��m¶թ��6Fw�7c\0b�t
�ο�ń�4�C����F^�������5�f�ĲuQ�IE���_�F+��F�ә{=�,�Ҷ�ע��:b#��<���&�'���a�#�FU�-�!VL�W��(/NTP�(����� ����wu
���9у/L� d��Ne;�!ť� \1��S6����,߱d=[s2��	�	/�W�Z�!�\[�j�-]�̃��t<����.�O��ؒ�����Plѧ�*%�h�id�Ǖ8D��g0t��)���d�������`�9`���E�pl������/{���DV�m鲥>�Ln?cc�6�d���Es���
�B6�Ц-0�N�W>.Ta�L	�t���(�'�vۣIVP�s�⎐N���Y�A�N��Xݓ����+u!GTz��Fe�n��4���M"B�����.��~XX�w8�o�D��9����w���{^ÇzD�b�������\���y]kGA�R��	r�	�ס:R
x�� 
 S���p����jVճ����o��=�P�m�>b�G��i�
��*�G������|Kqʛ�BVv;����$����iLi������u�o$'��%�<1��o��\����y��'-+����ױ�k�n���vZ��	(}�}�km��徙֮]�Ʀ���f��[�~��<-	�G6&�@�տqkK�D���f�p����v�
���`m���i���xq(����"�9"]0ޓ���y�qn�:���v��y�}����O�J�"�M�﨣��F��w�^��~�Cr��,?������sX��\s��7��M��W����_��_�b@���}��zPԮ!�Tɂ�����*�G������5RD��5�C�9+�	��O@�G]޴v��p��,�JF��9y�q���=mKl�r[Z���J��)����$���MO�j=�G=��b?�'Avj�Ɉ,��
�F�q�Y���>���m��?X��%Mf�_�'�hc��?Psh��j7��ױ�?��f7�VGI���s��n^��Wم���d�(�sءk�g��)�'�z�]w�u�%�41��o����o61�෽�mnݱX���/yIg5[S@uY�>_��~�~7!*7�xV��18�4|-v�K���������{ /�	9�����VR�o,�D�����:2	d����C� k-��ɉiMTp�D�Ku�ԴE��=^\$ŦGy�8< 	Ш���5����E����iT��?���(�����n�����.U2�%�Ջ��:5s��U���k�:L�\y�u���-�\��ǾZ��w�@~����,bE|�w��C=���_b�]�^�EJ�ܛo�E��=���v]�����l��n[~��=�ȝ�>�~ g�v��=`䙝Y��$�)u�[�f�x�Ŷ|�R�ԎO��&=�ӯ[Ln��I8�����#�����޸%R����]�S���?���`_��ל��~�Wx!1<	Tc1<R+ƓO>�/�>�����3���ҏ
����	��Q����+�O�����;����R��I ���תe���Tc6���j,��CQ����Vj/����}vֲ���l���:)q<��K(&��}}.*o)J�n���uia=�n��s��݉-��-�J:n~l�^_�)k�WD��9�6�VS���8i����������#��j����'�3��ח��d8��H���E��e�'�,Kط<�E/�K=`�r��V�q71:n�sn�'}�L=�ܳ������m��<kU:yy��zꙶ����C׮�+��F�=��;��IF���>�9��N��3N;���^{��Ǽ\0�T�+����\d*�L��)���,J��~�}��fk6�Q)���
�"I��Ijg�3Z��<�x�#6.n~6�m4Y�p�I�X,�o|cZ���
.��`��Nq�9)g%�}�"svr<���z�Q�����VI����}���I�ޣ3���l\��{t,�4~?�WJ�)�K�)��g�3������͘k�ǈ��ێ��Ȭs�w��y�������q��z������V��hbZ�d�o�fO<�m۲�1�ի��I'��%����)��d���a���g��c�G@{��V���\�d�Vl��ەW��IcjĞM����~b?�$ؓ�54�'|��m����9�BW e,e5ؖŀ�Ǌ�aA�z�E ��&j��I��5im�[^�="_XV�g�Q��6�P;:�Pu2p4�	ୈ�a��4��HG���y�+/A�wI��r(Ы2\ץ��=<)���p_L��1�O�ڪ���;h�e��[bj����b��mt���^�!Gk�!��������M�~��ݓ���^
ts�>^�k^�;��#lb|��Fw�/��~�������l	r&I����y�A;����QGW���w������.��|��>ϑκ�c�+u����Sq���g����u62�ê��my��$䟱�]f}G��� ��:"�w�����9�W��J������g�E��br�>��F����{�x���}���*���;�Y����k�+�$'a��6T�+6c���덂Q���*9��-��_��L�+����P�G���"��9aD�"���1^2�2���|�
�1��n���(���X]���2�w�����GM}�za�0x�r���w��&���3s���gG)q�?�"Y�q._����*▍���g�d)_�k�8��f N�y�+_�kO_y����?�coV�o�Ϳ�?��?񹈙����?:6l����Ϟ��H��#���Y�i�9�A�뮿�N=�,;�����Î�N8�6w��	!���;ow�!����j'�t����X5�?��F[�jȎ?�����4�c��J�W�1۾c��%�Ɗ�k�a"�ُ% ������C�1���C#0\�ˢo�34]��t�c�AZm']��Ϊ����<*���������Z�^fA�H����6��"]K�������X�y	��>/ap����e0ڨ�
}�=�s�;���E��k@��;�����;�)ԧ e��4's����#C�f�3	o�S�����\�����^c��#���:�,�����!u�t�MN � 6��u~�9�V�f?l�=ro�)[�n��?��F�G}O��Q����ϭ6<2a?���X�'�֭q"
��=�Yi�y�^��X��d��v�y��iR[^5���n�7��r[��{k���"ob�N�ɢ�8E�Jε���<xKa-�9����*ңW�EQ,7���p8a�ެ��Xp���ٽ�����}s�M0:��3����R@ΌH���Y݆�U��N�������)�/�P���ΊMlP�*��y��*�8��ň���ǡ��ӈ5�E��#�TВ�'�C��b{	�={�uf
 �N9[ڿ�S$�u�?�;�:����)��X�|'xM`�[�pσܗd�2[�z�M���FQ�u/�����a�Q�u�s���`��w�{lx���v���E�����w!\��g�ޘ��ݝ}�����NZ���`j4�=Ѣ\��-O=h#o��/��{׻��X�� Y X}�����z�j�k�GKMp��ǋ�'��%�c�_���V6�h�6#ŲS�+�+�!�XL���*�|����U�}a����0��RL���k�+Ll�Q�C
4�q%�s!.
���	�+r�9��I	h�u����B�뭲[�e{aÜ�q��}W_}�{��f���|�����ݣړ!�9�{��s�l������MM&�0>�{a��¬zg9���z��f��
�x¿xT{�����{��ղK�V��*�_�����¤���P�ȳ--���
�����eu���{�m_�e��K� "mADE�b�h���-&Q�����"��b�-�`��BD�FT�" ҋtv�������|��~�9��{������ܳ\�ַ>�yN���]�AY�x��%/	��������,���k��qՒQ�>N-��U.���f��Y�x-C�(N��9>�#_%��lk���bm�m��R�f}e=�l��g]D�)t��8�����|�]���g��X���/�:�|�Qh))JUH���<ήJz�ĸ�X��u v�׫�<某��c`YW��؅�[#��i�9~:xp�VdG�.}� �>�>ѧh>*l�e�;4`sk��q8�}����Ͻ�֮���2d���� ���zu)^���oV�':0X�n�`X�|��$�H1�É- �r����� �F-6��A�bn�\~�_X��$6�`}��Q֐�?Gǘ�^i�öYub[�2�═��Aơ8h 9.�Hʿ��|�X� (�FP�V��H|��{�j"��~А~���x���V����7|ܾ�8tͲB.tL�`g<LQ5�L��;5�,���h#[�<�s��ʿ���a��Yk�=eH���\�(��?�nr�c�Q�hw��.ŕyvg�5�7l�Du�n$���Y�/�"�����X��<�Jޑ�nl���۲�J�2�eO��)���wo���w�)ny6]�W�8�)���1�0��+R�ʩ�|�{ʽ)�#���I��O���]�7{�����E�Ѣ^5R7�L2X��e�s��$�|�IV���Qԋ�o�L{�4��e�����ްt�n�)8���kV?֬Ò�W�9�^����%�Cm�3<��6������������@ ^�e�h�Ǡ���/FȂV�2mi�T�b�J���bT�H@_!�H�Gh��RӾ&J|XM�Q�y�b�",�u���.�-PW�����`R����V=�Hx�I���Q9/���JX�t����[n�3t��y�Q�T��r�%��:�[�떱��X�^�[���7|���8&�tW�.�v�����~�oX*ЬZ��/n����Ï�vTN����7��Ƴ8w�q9}��3Xy�ќ�MqKK�e	ζ�egY��|$P���լ<��I��S��OsǗ�����>'*��������|�0��.�̌=��>��]tQd�6�o��݌qu���¦�=Hݑ��m Ϙ����;<�ȣ����]����"�2�z�O�4 |7��J�և��7G��~�3�mrg��w���M�{�N��`�5{n8ꨧ���=.,^�gN?@?OY���s����Y��E�j����7�y��=�4)ShK[���p����(#�Q�=��l�Դ--,�5����WD�8�a����m�<(�����%��P;$��u�3CT/a�=��fox������j�8��#�	+��:�ظ�u����?����R��"��dfZ��&an
��/*�+���85�}��ap�?�ߡa���	kW�
�7�7��yX򥳣'�^Eϓ*K�����0��2@��Q�*���}p{P�L�|M��a��2��4�k�TO��C�7����a�\���e3�o�6jz��Z���`�	ƭ�>V?�"���+W�Pm>�⇹_���I"�s�!����懧���s@��Ca�ڧ,��v�,�=�[�(���Y�B�7�䧡�ws�M�Im�����vا(��	�	��VC�˾���j�S��SN��˼��¬��aϐ��VK�x��|�;V��V���e��x��h�nv�@�ɏ~�c��a��Z�CP(�n��۲������M-��q}�-ʈ�K�N{�*�s�����{J��n��p�Yg����}�d��#�/E_@��
B'�+�/�z
�^t�������9+,�u�%�}�'�,�������_�첼��r$�-���E^�&���/̒QI5m���L����ζm蝑Z-�6eE_�r�e�a�k�+,_��W��>��O�M��T+�_��B��@��mT+����g>q�rN����ծ[���%�r���4�<��wɋhDR+	kO�,KO	6_il�`����%?��U�V@�?0ʒ�_.�x�ڟ���U��:0����y�v���(9��Q��Ch����E����?/��� ~��*DЧ0�{(���;�x���g��Hݠ}P��_�����|.�J�'�]ͳnf �:�R9>~�!�ED�o�`�P��}����eM��R��c}�N��4���~�㟲���^�|O��Ю���#��!%)k��MB��e,K��O�h\�"b��7�#̂��0�ꈕ�+6=d+
�}��TV�k�b-�����yN�f��G��U����
A���3���n+�&������O����?G_d�Ϫ�):��/���i2E�U��v�IR����i���f� �{O-"cf"�r�?�A]�=B�_��W�k����eFY�E�<?��,3\{�V�s��#?��T����f,�_�Ѷ����0��=���n��PTG���R��&��o��P7�6����yG��޻�W��+��s��i�Q��C�AT�°H	8 7S��$�E� ��J���ۙ%�dmx�6��-B@=�M~OG��X4"
�RĈ&����j�,OO�e�����h'���.ޞ"[���5LjI�GA����������&MGƃ����i���2N��E�k3kV�Q�Jɐ+i�r�r����W��($�y��mA96%w5�՜E0l��/�B�&�\��%�7���1�ph��~sK�H�:���>k�H>Č��j3�ᶞ��?U��9�����P����z:�j)q[�,�tp*$ �k�z�ue�{��&Fb�t��(�d7���<�y ��+�q�WGY�ry}�F��� =7�?��s��t��X��u�v�U#j
�� F�LDj���m�r����H,
o(t�SnO���UDcK�Y�'B҈:z2E���;�1����KII���@eT�o�q$�~�9�OCh5Q�0�<�@��H��QJ�s�/H�[� ���/�c�h/U�(s����z���������>���)���
���>M8;\Q�&WR�,��lT϶�,�� �b���k!�|�;��c-fċ��ѷ����',E��1���[�Z�|!J���X�s.B�t=4h�Y�:&Ÿ5���h��=T�������Gu�X�;���Sr���)���=S�xD�!�U�Y�IcE`_M>٢1�á$;���б+��ΈC��ԒQ�D��'��W�u�Um��)<�n~1��8 y�˅�Ȱ5��f�%BX%#�K�~���=X�J
�n��M��Dj��V�K�����?KWm�MT6��ь��U]����\��)�	�w�+m͗)�Q4ΙE^�p˾� �$at�W�}*iE�h{���qkI=e"��m&
/�2%�\��EMqT�Y+�;�[�PQ�Mݴ��L�z(sQR+�9ޘ��-诮k�/�m1f+�w���dS6{oᘸ�,TB� >�篙Oו,�&o��y�	�Q(��s��)�Сs�O�_����2gNOn�#D4��Bm7k#y4XN�Q�/��C�1�a�V�6h��e_�J=�7��Zr1�0)%P+��>?���)�jV�7W7��7V�Z�u����4T���|����{�M��=��1��n6�=)"OC�WT�Ÿ���0��l-�E*/�,�re�v�0٬ �os��$����>,�d<��Aw����U�E/�!�@��C��X ���/}I�m��ro��]}��Vs���dJ=��Ʈ���/�xw�dd�"R� �'bl���$2BX��x��DSH/��-�7.�o{z�,�P�s�m�W�(�]�R��!:�d�y%M�p�J�J0d��\�aK�A�����~�s��y=���<�տ�Y����@۰c��3���Ot	B<Ǹ$�c��p��Q����b�����n��-��1�T4��șlM�k�B8�evi�x|�+��T��RMR�w���B�#d��q�$�uHť�b}�"�h���Ȫ'�@� cJ�ʾA���d��>~��*̼�9����5�8���d+���IG�*�5�&���Ƣ΅��k1�$�ܟGQ|��������x�5؂8,�Kc0����馪[ �a�m
LʉU�1G;;���\(��P�\�|LZ���u�!�ƿ���Q)���l
AC��\JW쁡T)��;�)r�W.���(&��A��H�=�C���{p4����h������g<>��̍�&��8Z� P��j��eU�I�s
x9��;��H���9)t)r>�&�硲*���#
=�O���X�"ߏ���T�E&[��ĸ�CD��*��h�Z��
z��-T�̪/%#�Gڽ� 3J5����ǩ=V	��~��&��[����\�W�Q�y������5)Z��������aJ�T����E8��Uμkiv���~���7�@�����J��9�ƴ;�o+2��x�::+Yf�ìl� pߌ�;k� 7Tqq���F��7B?�Z#񿑞�ږb�����|%<^��5�h �M*���B�c�R��������H��EM��\�{�"�7����;�;O���;�֌R:;���x�o��!����iҎ����g�C���Pv�Vݛ��g���c��E�wnM�y0�chA�}�g&�����3W�N���ם����`�ީea+Bf�yXI5A}}t��2�s<a�i�����z�IM�3���L)[��m�H�T�)e0�5��"@
E�SL�m�_�BXF%�)�k�c��L��SD~x��d'���O�z�a���m"��V�7c�X�_罴����}K��z'��|��exoK�TA��[�mlb�ް��'=J�x�޷���ֽ�tY�=5��\�3�֊�(?'u���|�ӣ������ȡ�S��Q��T�F������Z�q�CU�$��y�Y3iy�!����o��Ψ����)nx޼���a�:KΤ��(aҹ����M��h�7JVB,������ ��/Z�>f_T�� ��%哽�8�9mmry[$O��J9W�G��U�x��=�x��<9-�x
1�Z��S�L�xX�{=�Z��S��)q�v��&)�V�I����"Aj�a���[�$)%�v��a���c�h1U�I�� 2\��&��h�VO�q�Q����PV璵��r��y����s-,M(��`s�V����:`�A�����,�ߕ�����p�QG��sS8]�\J�}~}˯��<��Us"J@M�y��3��{��lq Aʊ��_n0Pߔ��58<���@�b_֢�W96S`�|����~���� te�q}szYt�WŅu��3���
!�d���������d���־��V�1�R��� �c?��f�7���crkI��b���?����j�	��� �[��ih�/������B�Y/*����ہh��K)�)��;��}�1F�ĢE�æMBGg�l�y����52+J�X�K��a��/^b<�rw�m�d�v�a�����y�T�9�~��������o;��W�J��q���w���ۢ�"��|ޚ�R����)Z��f��Dy���yL�"�u�$W�����.Y��&�S<~"��H�z�/U���@D?,�e����{P��M��D����8/�4�y`��+�YN�o-��A��-��Uua7�l���x}QS�1T�e���3�����~�Zu+�
�y���c�1Ѐ�)��y�q����~��[r��$U/'�iXq�I3��Be�%K��A� ���AR��eɀ%{W�^c݆@[tvw�=�\�X�$�_0�������������{��^'�/pMn��_�j���Q"�R���/���(���b���=yWq���B�ޢ-�#��믿>�
����B0���U���+o#���xg��Gl�	��ҡb\�;�L��E��Uա��>g�y�s��1�W���>�_g�>���=��¶���q��?�����=蛡t J�����'>�<Q�y�E(���;#r���[��H�QI�D�澰ے]ü�¢Ż�����ʹw���R��k��^������J�ț^��4gx�s�-�y�TNK�~�âӢ��O{z�k�ea���V���f��C�A��.}<�ce��DV���6@��XZE_T~>\����mg�Z����?�c�¾Ta-*
�;-@=	r�P���*>?��#I4&fb��6�B�\���?F=lUU�f[%��,a τ���%����w-(|?��s�T�2?-����u��`h�m?~_%�Ѝ�������*��g?ks�¿׾���P�P?|򓟴�#T�ƴy<���#?�@'��=em��֭��"�i���Jٶɼ��l�΄�ǳ�O{��L�ɝ�g\�l�p�����&�|�/¯o��ݐY�������=�����p��Ǆ�p��X �|�t�bWEA�k���lٲ|" �JV�౎���'��mU�H�6����,l!���F��b�ɡ��呕�a��}�"=��������~-�o��|��0ط9��prȰ��Hj!-yL!��rHߏvr�c���g�����և/~����LY11��ΒmC���ů;���SO��:8���^���/��b[���7m;�9A�������@�>��G�7�����'���=��~����"�(�:!�C����|{z�V�a3^�w���`�شV���n��e(*�êU����-���a��e��]�f]�ߟ�8�\�.�}�����'[G/�w`аYYY����c� c(yؖ�+R��OwԶ�jR�*#�oB��;�p��z*�4�)������p%+�V�U#�z)q��0̖����]��C��ې0�1E8������'yY\~�������ֳ#�0.ޠ8���z�E
LCu0��ۻ�=��*�a�����Ɯ���S�ׇ˿�p�	��7d�'�n���p�]wY$b[��i���&E^p�E݃��|�����/¼��a߽w���#a��}��b��֮[���p�?	���ߔ; �fbrr� u#�+ĀO�]A�����}�(i+�)-�e���"�C�������~7S�s�N�<GOs`CV��5� �~��hd%��Y��?I�Y�U[J�Bt�kr/��HG;�C�����cm���߹"�wιa����&Z�ᔓ�̛֬~*=�x�4*UxҊ������Q�$�a��Y��:�?@+�p��>�W?�fU�я�.�=��2�p���L{�J�#~��K��i�{`s_�;�ۚ*<�όx~ظ�'fq�rW6[l���u�6G��Gm�?�\A|��Y�SLX�
��'b5!�|�H[��-�l��hY�SY��y� ��X�a�0�ը���8��Ba%��b)U�fϙ�'�ߓ~/.���^EV�x�V@�/�
�^w�u����N���뫮���,���^>���Q � @��#�S.U��o�i�c�°�^KB��ު1 ���\w��`X�p~����-w�{����@B�ΪUOm�M{�_
�M��;��sٞH�C�#��0��qY�������\�a[X�<'	,�/��~�����;��=��!1��f1`��җ�d��3�I�D�ôe��p�J��h��^1׎DB5�bHJJ9�laӭtf�
��BZJ-yC1Z�n� �؜ΰ��Ѝ�T��I� ã�?���B<��Wq!�hFZ���O��-���7�l�n�Wy�w2�V�ZV=�xX�����t��l������T�2n�Zm�E@����L/�0����c�3Ꙕ��p�7K����ņu�CgY��MiqqʤV�6��$q�2B����� |F#x��|�.����t5e����
�Lm�W}�#CuYM�=�C<��"�r�`dl4./�åa�XH͈ޔ�5\F\ �� �M
?QØ�@�P�ƅa|��;�y^�2��z����s�����/��'�c��) Taz�CwO�u�d΍%�nI�4�
�Sփv�k�L���o&)?�4������Z���S���:-�M���v�OWGw�<0��ss�ӀQӖ����4/ݼ�+�s�9���~`�_����芧��֖����K�no�<�4�b����Q��r<�h�1��D�G?6[�5*�ٶ��u;O2�>)e��Z�	`��::��M�_砤����@;���Ë��E���/�x��q$��k���4�+c �Q��e �}�O<�.�E�ڊ�Aӿ�=��Pn�R����`G+{����ʺ6̟7� Vs,�?��tǬ8@;�������M�;��I� �"�Í�"O��$�2 (���#�?���?��?�/|����W��/(���-����S��{�.���6<)Z�C����V��k�eo��������'�������2ۢ�j��;j/(+%��E��*tQ�y���z.�����WCw>#�G���X?ߡ0�a�
ݺ��tu϶�J�fx�����5{j����ua�^;�6�gI���%�R���C女p���+��nV)u�q�psX�vSXs�TI����6�n��=b7�?�b�<n��ִR����t���Ȩ�;�n�.��_�o�}�C��N+\$���e�cnˎ�ɄZ'�TQ���(i��0	�t'�P����ڐ%q��*Y��?�i��xF���O	��`t!�d@���.� Ý$Y�_=Ҝ��-�fT�:�֦�����a}X�~]� \�g����x��C��Y��N4 ���MF�F����	�6�
�V�����{-�#���;�7���W�5�����Īա��k���ƀ�����B[�]K�i��s��VD���p�aO��zsX�a��*����[騄����~����ͻ��s�N$ox�����jx �@l����g�"�EEBB���Ԗ����5/یs�_u���������uM��RW��U�P5mi���j�����\��_���Z�v���-�V�%�<1�j�ق�!v�����I�U��9�<]�O�����{�Wx�oSX�iM6�g���U�[I�ݬ�粽�I���Z>�߰1�u�=F):���d�S�eȚ>몃�?�C³�����Ǎ��'J����3kd8����Z��QO;&�Ǟ����k�F����mA�g=�n����j� H�PZ~���t����-h�Xpmi˶�o���� ��w������y}���z���ʯ���Q;{�_�|��&(o�=*��>�ݴ�8��_g��W(��ܠR��\H��/|���^�2��R�c]�$1��0�|�~��������t���/<����xU2~��v[N{�s��
s�.�c�����]w�6�t��;c��5���T��!�w�WZL~Y\�I�{���|�>�Ʀ��G2g��ea>���ub ��e�p�~���VOa��
�ָ}(�W���:5ߞ�(�����J_O�M7�d�1ա����(��� ���O�H� Ҿ���U��J�����i��R�导� ��9�=�г�q�f�!`���A�0���9>u���W_}u�m�Ea�ys��y���f͞V�z2��m�r���|�5����7��^{ì�9���U���o&iB'����������a�����a��9T�����oF��~�j��FTra@��+v��;��U�<h-�do[vv���
w�[U���o����r����zܨ��0~r�?U��ߛ]�z3�f����z�*�J[7��,���
�b���׿��]�O����(~y@ZL��^~��-�=k^\ ������@�ي�2cq���QGt�u��{��U+-<T�3��m���q���Zޘ�%��/~�?����7�����q��W��6���ׄ��+�巈���������fx���;�>������28���w;�Iy[ڲ�ģ{<���jCi�ݼӮ����m�$���y��6��gaTY\
`Ͱ��l;�W!��"�c~����I'�d�Y��	�b�Q�N��������O<eq'|�;��:t�;(b�i����On��y����S��*�^�7+�R���m��fϝg�W^n�����u���LY6i��?��n�:(-'��!]$�����>����f�q �/\`!{�ψ~�c3,0a _�5=`۲}e���L(��̘������@�u�E��8\�`��vBj�S�UΊW;�ݲc2�Y��r�c�D2t-~��`��>I���_���l���MA'9�o|�F��^Q徘z�B����|�*�n8萃��˖[�?�G'<��#�E`4��\�6ܗ�3�B 0s;y5asey�jg�ǒ������X7��?�x6,2���B�=����W�j�\F�O����
�����G\�mi��*��0��ϕ���	[�V����%�����{.F���O�f��Y�[��A�VT��OA�5x.�³4jBA���O�~�к�{�F� �
���Y���Z����O�G{4k��:+{h�����z���xB�X��}��]�5�`-tf�a�q�ש�Q�d
��J�!i�!�Ց���^X��/�� $9������e��V��(`[L�V�}�X�FZ��w~K�@�������	g!�<��/�	���5�暩�����:�*�B*���{�"X`% ���~};P��HH�}�mn{J����3�Z�V���Xv���ζR��Ŏ�ي%tS��
QV�(�T�b�'�ݡLq��ϊ���H�ߏ�C�{�Ï~�#�ü'����J~r�$����c�CF]�і��7��V�e��vU�F_�P��J�⌝�ʟ�݄m�TMNu�g�k�E�Ɓj^,}�9��L>�z�<H� ���FZ����7�).&c	�X�WyAS]�#XQ"Ucb�
y�y����C��Ct���#�+.�;)�c�>����[�o�_�}*Y�R�o���']F���X�ԓRP� ��^��͏J�¼s�k&�jod �����_�����Ð�}��`��<PO~+䞌�����1�כ�(���?.���Qyc��^ײ�6�^:9�܅b�@�(�z�[�j. �[�����e kLx`�f���N-uo(k/5nbK-�$�G�=��A�K��N�Q��{:�f�Ų�EQߓ�>
j½p�[XB��Z�@-�gX���u����MI���/�B��g����D�@��(} �]�V��9
�3���[���;��1���p4t�J6�E��E#��5��(es"d��>q�_#��j_�̜a�R���w�{T�W�͇?�a3�t}8jd���Y]-;���%���]u��M���p��W�(� ��|��A�í�x}(��hpȂm������0�({�Ϛ*�r�?�V�T/2S�FEp(D�b��𚸈��=^�Π��E��<(zAh�e�6F)�d|�����I����ڱ�A�����D�_�GJʟ��$eP��@%>(�8I��WD��͵���ͱO��fVO��V�Ŗ�R�fd�o�3�<7]SY����~�%�Y#�Zy`<��m��fc�^��k�u� MhgFf��yK��rke�+�Z��/^�r�/p��`<��ۥp�&D�%$&?�#�`��R@^���5�e�*l#��lb���>�*�U�Vc��-�֥ב��B�d��R<\JQ������^�F~�����Pl&/y##0�P��țsF�)l%Ũb*?~�@d���K�Y�v���&��l��ª����Q�@�t�t�b��+Ua������Gख़��gˀVV��f4��6���暊��z���sm��3����tq��W����V�~������R����uq6?��=��?�IG�&-����($��m6)E'%���>�z�>�.Z1�k��&G&�X�:�֑Gi
��@��>���}�/�]�\�ue1s��7�Z>���H����
e"�N�FU���0$����jH�Q��������1L��������<\�7m���I+��c�!/Y��pH�o���?��&a;o4H�3��a~�9�;ƒ�����FyzJ��#-*�Qa��s�O2q�~��W�IǺ�z/r~c�(H�,�}�))�)��G!yإ�<gx+�_�c�X0��؄��,�~eD��M�䔬���I�s\�dI�O�gAn��Ip>'�A�)�t=��gk������,�f��ZȔpTX��%�s���t�:�9'�!#�EC��z�#�����M�K?#�~�;JF�2589�]���,5lJY���Y�w���04�.�T��0����tTlQiz�uBz���jg�j���9���t�VR�Q��ku��ʴW���8�}�Qc}�V�����z)g%"�KO�UB���C�DV"x��+7����?
DI-����1��krj�q�b3-R��z�rC��5cA=K�ԑ͔��x:&ŏ9V�[H$��PD
1�D6��;j(�筧�{�~GAWh��=��A#��b]K���Q��(�;�<�&���`S�V�J�S�HcEH1�-���܄�Ac��W3=�~kԱ��fe�Q{���к�J3�߬·R�j8�a��ڪZ�IȔ��:-'O-B�db�zG�k�'��/�������ڷ��5����J $q$pa3��w��h��0)�=��::Owg���j�����5l�^i������2���#-*����^�h�q_�&���r�0���=e�g�CǪ�i���PЊ�9��E��YH�63^�o�;
����N��!;ϸpu���?d�,�t)�Q����@H�{�+]'��3؊95��0VA&Ǖ�sOZxձ/�0�E�;�.�nʍCc
�:�s�OǤ�u4�Oc��i���a�&�c��]w5*VU�z��Q�d78M�=Q�����h&��w���o�a��e��
ӣo�(�&�b�<� դUa����)�YY8R�,��$��ީ�gx,�����'/O�s&�
�
!�R&��QQ�����ߔ���(�z����^�+��<�Ƃ��p��<U�1�h|)�%e��������RE�'#�X��?�C���?olճ�uZ���e�]L���	՟�Z�9�:�����PP�'�Y{�4��	a�Y�������?�䨄>Jm�:ʝ��m7?���OJ��P�E���_V�x�]`�KC(�j۷y �}Κ+� �u)b �� �_~y>0&�:�.�&.�L���g6Pe�kA�v���,]���j�l����W������=TL�
�M�ܟJ�'�T�7�wW3"��b�0c�q�x� Y�Eԙ�c�#)�E~"D	LY���9yT�Dqr���sնx�׻���TG)�V��/��\�Ej�:�K.&x՛�!5M<G
�)�$���+�cW��y�ᤓV�=��==�J�7�m��Px�Ǭ����z�Ø�[XX�ɴW����]mC��3�8I����n����M�q5N3�==i,��U�BϬ��Y0���B~<�I�l 3�T ��&���Am1L\���Kp�f	[m_1��!��������O����b�^� �$��$/�Rca*����(�K�$����Q���E�(�F���R�0�S߂r�a(D! ~ON��2d���z�������﫝sJ�Y��XT���t����W�e1���{x�P��T���q���q$I��!r%[�jIX�d���z�<��p��ׇ+���NW7׫�<i���6��M���I$��N%��o�J]�d
��|����c��@�%�l�ޡo0~?��B�pË��v����D�&�?� Y%*�A��'� ��K���	ca���<|t��欣����u��ӻ�
oy�xkE@�[T� �(j��7����t|��b"EJU�A��X���D�U9	��(��Έ3�3�󂹧0k��TU,�w�qǍ���ʯ+4+��T��74&tnԃ��cn��؇�FOPV�+����ܳ�	'�8!�KI�˥Z��;�d|��q� �6�<�0�<��ʧV�cc[e(�ZCӗ��l	��>��/�ma��w�yG���_��}40�
;����V���?�~'R'7����&�,f�;�!�� 4lrtt�A�i�X"�e�w�.U�
��f�2�����lU�����
1�z
��(>�������M��SY�:&�z�F��>Wa+�����1I�,��_���S&�x!�B�SS�õ������4��&�����3��R��������[��ݏ?.|>��`���o��d�bU��v�iv�4����(s�'�|bڏ ����3���w�֬[�ſ|��ê'�O{�3�ҥ�����-^�]���Ӱnh��e�Z�%cc[�|�֝^�����љ��
+W=���DK�?t�l�bQG�7�p����Uk�QO?6��*�R����N-�<
Y�~Mz�bXF`�{sT���#耱EO�J�AU����G;,|�<����ĳ��8��"R��{x��d�VP�����E���d��ZBQk��W��ZBaފU�x�V�.��'�=m��&�E�|\��Y�F��ys�KKR/�m�������4W��|������}O���Ҽ	����V\��`Q�oi�R����/�{��a]T��w���9,�M}����~���p֙���S�@����([�ʴW��	@1���Ι3;U{�o��M��H�Kw�����?�)~��.�����}���?��!y��7c���z�^hȋO�y6YXF>��cͶ���#4�X4X��,⛅��
p�F�E*O�;ؤ�*\�7��d�Bl���a��yy��M+�UQ�D���J�
�H����"b!-g̞�{�y�Ɵ �����֬��p�C�5��r�~<�Z>^}������o��C�f_��O��p��[N�s�?�lI����
룞Y����_�bx�E�	wYl��#;2<�Уa<-�g���	tW��K���m
s�v�[n�U8���򽉟�5k��;	����as���zVX�nc�����z4�<� m!�x�	<4yx�^`�#{�'�MdYy���������O����C 5Ƚ2���h�d����^���tN�!:��]�"_Q1Vު�ڑ�$�����mC�WJ�U�L3�7�"2�\|ިH���0��[woC�	��d[9~�ܥ�{�dk���И���?�"�EO��^t���1�c98�F�0�U�m֪᷿�9��	a���>4d���ӈ���V�z<>�V>��z�r곭Q�A~�ӛ��F��Z�.ȴW�I#��RͲ�W���3<�أ)�H�ue-�Y��G��ąN�E �o����`g�y���TSx�'���/�5�җ�4��_�e���'ێ�j)�V�r�-,N��aq��M=�d[�SY|�{�e��D��?��Qdx����˛$L���ӱN� y���i�B����~���r�O<�8��
�%��@�+W��{�p��ˣ�9/.��3�� J�[�TaRl�J��<��,���.��#�?��p+���W���PO�B�ء,�����!+��������>��+Z!�ërχ|'�/I,P
,x~G�׿��f	(^���b���M�����+c���V8g\e�QԬF��9��'ק��L�թ��D�PR
��o�C���y
)��~����/.J��0�"O�WI+<Hn���%��+����}���Q�j�ĸ�GT��
�R�3�W:�EtpB�8�fu�����A�E���<�#�^����jQV�j�u��7����՟X�]�ܙ%]C�����qM�:�8�,wA=>a���ĘZ���7B�8U*�jB�4�!w+�˒Ŝ#�gC6�ERS=��E
��'baf,���~�|�m��62
�Qb#�0��&Y���IǦ� ���檼`<\B?��Q���+�'�=x-�a����\\l���e���`^w�Q���OL�uk���W��ು�ƥ����[ݳ���`�YJ%�!�^*u�M*UR^n"�{!atS�^���O��2�L�>�{���y��U�F�8�BGE�f�E���L�\�ĥ3�K^���O~Ұ� '�˼=e�A߶�GDʟP�^O���Cё����~fFA��B񵒱�C@�`
���G�&��	'�`s[ʜE�ӷ�������T�������ƅ�V6�r�_�V`��j�~{��.:�3�#
�&���L�z&}�tRp�kf�ww͊�¡��Fk}m�Y��h�f�QBgX�;�Ǯ�W���?�'}�Ї>d�>&(�?x j�۫ց�(�y*%�&+b4T!�K�[U�;j�E�����F��-*��)  �G90U$���J�W�J�z��b�Ó��]:v��!� ����Kx�0F�(:'e����9�ȧ���k��5���:u�9���u����-�bŊlA������UO�L3���	�j��O��]ʉ�3���{Pxr�C��G�aH��*�P����[������ ���Zgq�f�q��)��(8٧>��N)@�>	5��2��l'%(�O�xK��
�R[;�0QhB2�^�>�-��4��c,����\�\�o��2�h�񊮗�E4J���Q�V�}��P��u��4�p��>���'<��á .��]�E	�gO���ݢ�K�,��E��v0b^H��<M9"�T�_ٴW����#��}�s^�={��5�+,�.�~���~���Ҙyq�8���1ǝ:����V�V���
_��YU	"ڽa񫠊���<jH��2A�Of�_��2�t�bX�8����w�(�;��d�c�|��4变r���ɂ��fAP������@�I�&���������������}����k3 i;��cC�^{Z���ݖ��_���0ؿٸ�6m���ts�qǞ�v�3��p��	�@J��3*�g.�O�2��:+�B��������0{ޢ��!G�E��m�;V\n�.w5���h�@�I%7���d ��ӟ��n�����  ~� Ą(E�KJ����SF䕨���b�0����D������־�4�CV�����lq��
������A�|�q��L���D�w���	>=���¼{e��KϷ@�v���s��>Av��n
#z�~���1��%���·{ "��>!���Q�0>��������]w�i�Ϳ��?��N�,�T�` 1�1��$�İ/`�%M���G��M�
!�k�C�3�f|݊���wb��Sqt�d��zvO�O�����X��w��k�i�j�A%��aNT��.�?�x��E�=w���:��|�!)d��6n�W�ϕ�_c��]��{+3��O����K�f4��=[��Z3����h�����E�ȨU5��j�0�:���M�!\pAx��^��o�&\q��k_��YLLmW1Q�&k�S�>b�����K�"��k&n9^xb�hdbiۂ��կ!��j���I�ce��NQ��s£)�*�@�d#��+�b��c���$�}G�yOD��"+��'���WwM�P�B��E�+��B�B/�h��_�<�����@B8��������E�r�,
R�x�į/�����;�1�c����)��H�D�9�1����s���crO�f��o��`*����d�׊sa?P��M����4��/_ȋQ�󊗽܎o�Ż�9s���?$<s�)mC��>�9�P� І�%���)4�zjB)#�O�z֩,J�:_է�7��$(�!_@�]Y)bGT�NJ�6��`�Il����@r���>` ��\��p�r����0Y�-�˕U�;߃�.J��	Cų��H������{r�RZ:�S�B�Hd=QX��/R�οނQ�.�G�����ENVe=���}�zh��q0V�@*���+�}��Z�@,[�0�}�7�*c���£�������LfOx�P|��zECq�T�KIm�k�����~��_<�@;g#|G�~�Be��wA{H���CW�f�q.ox��E�C,<���/�\�1(P� ��K�~��~z8ꨣ�;Jx~)^3���/䞆�Ȍ%v�����WX��z�M7�
#i<ł��Z!��TYV�D����o?+�Fi��]v�e�\�w���h'E�+\�5�Ӕ2�I�q�9�+_��m˔t�:�!0�Aqބ��;����;L���t0�\�Rǣ�g�{˓�c����(���̹�]����X���z0Cmϓ�),e�C2��T u���gE��!U\ �u(�(�;�qSj-����3�Q��\s���/Xؾ�	�
�"�f������?�+Xy8@�Qp֭���	�O���Y �sl?ߕ{�x�o����g���O�$�'bM�}��,,X�Z��6�	p��싱��x���x򋱮�t��w,:��X���g�5C�Z��`�q=�y��F��Ɍ�zZ�Dq�
kEn�o�"�M��h���{��)��b|>
�N�@�L�`Q��m-��@�M���w�-&���x�O~�܂`���/�{�7V>��$

YҜ��d�� N��eeyŞW �}Ja).�܃����X����+9=�2Tx̋�ڢR��)T��o��d�_�t>~�-��Ň�t>�影Qצ�IP¬�Q��΢ �C]W�	{0�x-CB�E�Oޯ���<y}�7�a#o��Ʊ�m��x��[����2�ѥ������m�$�6ʱ��x ��?����{��^{�:�	�1�(��A�����9�ЖI����3~�G��c�'���C�EI=]\YA
mx������c4W	J���X�X*��b�a��O֤� S[;3�G�_)|3�'��%��%7ٷ{�y��XM����x��5X��GǨ��rqY[���4pM��G�z���U�P�6R�XO�c��ݓ+(�O��ׄ�qY�+�~�H<��,:)1�g���|2��̞~z,eQ�#��Z�-�~z����w��[�K
VcH��C�}���3�SCH��@ʠ�exCL9,>c�1t�����Ka�H}��G�t���9/�/0w��_��WٱC�v����X5�}N�/�X�bDe[\C�O��P�)%��6�><���ذO�q���|#����nAt�"�|q�@#%��.��P��J�MF�Y�?ɋ�d�MB���)��OhY%rk-ќQ:�[ ��z�%�BԾ��P-Z]�da!����?�SM���J����$X9f�l�� ���D0� ��x+�uU��{����Qܗ����a����l�+FΟI�dS�h��'Q�,��(/ΗEoO�J�EPJSR/���ל}���kxl��d趾��ay�׍k�}��5��uQ�����cD6�[J����!$��'�M
�Ѥh�țf�a5��߶��·	������K1yY�7�ٟ���;�7\3§�w>������w�Q��uև�Y�Q�Ωt�s�y7{�\�� �cp6�z��a�&��\`o�!B�ԋ��X�B<�#�G��� D���`>~�d�,���QP�E
PP7<�I>a+/AJD������}�Rg�qFn��!��J�Q���cb`��!�K����-������^JL��(Y�LL��e>���d��Zם�1�u�@��mOׁk&��~�m���|�3��/6����d
�Ca��C�0Iz^{@?�|���X
�#�|e�)<H�k�H8��
s� ���J����'��SO=�ƙ��
E�K��s���k���4�4�=�*���xd�(SZ�8O�����d�)��v�NT��%ijOpj��a�>8G��]�앰ւ�ךk���n@縵R��8�������U6�����2R�>��x���b� �()[M\�A9�*B2%KE�X�P���ؒU?9�ө���R*��� U3���ۿ5�Id�*�^�W���T��hC	̕���Q����(��4[�t<��|�+��ҹj��9�""h2E��#�J�^0J��9�z�ߏMY��������gD^'���'>a'��v�(k�G��vAa�X\r�%f�{�[�iy��7���"��BCR��X�}D<�Ya%b�,:��\�����{!EM��d29��H$�-��_�a'?������Y����Lsр&~��镧���y<dybrJ��5p������Ʊ�� ���#���N����{�]w�n�_ F�m�]n�$��R��`��*(~Vᕼ�}�3dぞ�J�+�Ȃ�� ��N*�=�n���9:�f��q~��"�?�S�I���V:V-��/�5�����%��-�j^���,s�÷��"� ��R�4%�j[v�裏��|��W�DM�g'�t���p�KɃ� D �������*�$i+�F2�y%wQt,v����{����o�KȊW�/��bJ� ϕx4��%����Dj#�6��^"�<���#EĘ�e�����'j��v)��\�;�5�\����CM�Da�Md��Z݊댧���
eP��"IG|]�p��y�"l�U)�c[�7ҙ�������X�BQ���R	b[�����A
�)�%�4��fA:6���Ci�UO��	��|�BB�7�Rj�����
�u�%n694h}�M�6�+��F������*�qP�O�KK�3�U-�_�1S�L��>mIe[c�8v�R%����ڗ{�g(
�~*[A�YӢJy���C@��e��Q6�3l,��k��������ߓ��WS��Nŏ$�����Ҵ7�(V-1H�C��U�XWL\�4)���~�����b�m����ZX�@�����(�w��?�m�Qm��(Y�L���,��s�U�3�����a@���E��1���Çu�:>�x�0�_,����\xα���y����D=T�T�i���{�_� T�3������^n�{_4�s�Ө}���Ry0�<N;�ܪ�ّE���J㷼�-�}�z�8�[��m�6Q�{"�` ����+_�J��!�O|߃�(���/�+����R����B-�����q��m`xlM/�F�P�^��TV�ȴW��=�o�!g�D�z�*��!FK�"b����CDV��T2�Α�,�?������\�h<��x-cS[ƖV8{Z:�H�׼�5�ȧ��<�*h՗ZL�(�������s��/��3Qt��G�ÃT�f�*�Y��yHo#)r yU������/	Q��2�?@'�����d�Ax�5��0�ô�s	���	5�:���B{��G!(�6؟&ߨ������6�,��a���>=����d�����o_�p͵�U�O�tWg�q������MZr ����+?&D�i��&؃���[[W�R����B��b4<h|M~������X2�Ǌ_(���
K�"����`�\��j[������(�ָ}Cx�����k�r�=N��y b�_08Ny�~�C'|~�G��A�!Z T9��=��XX�,>$�	E��R����G���������Sjܔ��Tf��/%;�寄����!zx%!b��Jx�b?ȥT��e���-�&�`z��9���"���B�!o����G����.E1���6a�f���bbX���)���R��<Q��W%F��4O��b&���������o��
ay"E_��{,���C*�!���������X����u�[��Vر�xE�%�N+�B�o�<�?F`؉E�@�T��^
����ʁ+�䘚ë+������9dWPȂb����rDC��[c�f��I��}c�q�>o��V;z��H�n7�0��m$�ے���3x. H��o�h�IE�+���}�E�����ٶZ�"���V�%�g�D���E��_�%j\� 
���k^͇<���rQ����+�s�8�����M\vV�ǟ���ʿh��l7Ӈh'[!,!^snX_|���'�{<N�X���˲?��g���|vu�\G�F�o�zƭSA�=�xA6Fs��E���7��DSma�;�!h&r�Ց�S;p}��s�?�g[R�u��1(G�X��ͮ� �,�,�(Y�� �4��<+�((*�����18 ��,�Z %�C~�Lh��&d�3���2ɇ)?��T���(�ڷ���ۙ%���TM{��lugV���n�s)��9_Q�X'
Z�Lաk�I
���iʚm͝=ǬtQ8�j:=�����r�-��ũ�dR<ZU���X�g�u�uR"�� ~x��!�Z�#+�,Ă*ب�rK�E`��/Xo�Ḋ���U�3ް�?��O�7�����_��_�؅�����YX�4Ua|���4�-�U^$h1�Gq4)���2��1I:�!��7F�ƫX8U�"�-Q��z�m≰�����_)猻;��k�TJ����������Q|��^���M_��}�K�o\V\]�$s�`�z��>���d��
b)
��@Lo��f��O,�F�����!V��a7�/y[=g�IQ�y=�>��R�x��IֻN��#Dm�X��(.:tѪ%���7�$���XM�W�1n̂��@�?1��lC�Xǀ�[�2�+'����u��	H&���DH�?IGwG��ŴW�q�k��������I%����'��-Z�>���dՖ��N%ٔ�U��1}�6D��Ќ�5�W��U�Țc1�dl$�0<��9�Q��W�V�~݄�����L�o$j��ppO�N�?��8��҇�9�I��C��#���F�TM�Xt�z̿��=�� lKy.O�k�&C�J�<Ť�3��.�b�?�fo�K�B.�X�r�5i4@}`O���C���)���7�֢��M����ĵ���\CV�g�(�3AU��X�R^����D�阽���,E˾���S�Һb2k��ux�8�h���W�D�"P�9�43 CUOy �k�Lݷ<�ƷBA2<|����YO���VD��+#�-wf�T��==s���ٴW��Ty�[�^	*�3�E3$#�gE.M�9����D�)�llk�%!�����xeQ��E֥�s��e�Y~!Cl���6��˛%�&�/
�
����+<!k��J����\C*TI(*	�1#��S��s~?���י�&	UOR���:��"f�b=�>�\�:O�_a��G��O+���U;Ey�y&zD����n ���$��Z��K#�?U��E4n��"���_{?G4�$;��/gƛBV�����{.YR� �ښod�����7͟?��M�Ԓdf��+��H�Q���׾6\t�E�$D��r~��sP <�LEbp���z��$�'��T����b"���7��h9u@Sӟ��!�g�#��8F���Y��9%�E�,�&�4�t}�U�:MT��<:mp�����\�׽�u6>�؅n^���ã�?6�8i�։<o�5����ق�n�=������O��{�d�ƍ��w�&�T���D�&%���Lpoa1�9a���Ț���@�(!rI��	���g��_�z����R)ԉTVń�Be`�9,y.$79~�!�bƱ�:Y!���3Q�L�+��W��ն/q�����h� ����7j���˾�e�m�ehK#Q"]p�Y�O~��+��v�+���-��Z�7^�C�"k˶��1`���y�ؼ����b��C��v)U�i17�p���k� CNm�JHM,A'�'�^��c�'�������
˱ `q�|W��^��(�a����J"��K/5���������}�5�� ��7����>6�����!�EcY9�ٳf�{��'�-Ӟ�����O��v�i���\��5ض�'f[FD�F5�'!t��=R�R������ʿ��  �IDATK|<_}x��Ǫ�E����C$F[BO�ࡒ%EZc�&�΢0�^Z�|�J�m�d	��ZQ��9��0|��9F��.��2k���9v ���+̪�C߄�[{N�.�gK�-���u�p��ϸ�W}��o���GN?���]u��/]�p��(+� �k˶��v�!t���A��4)N�EL��_Oi��P%�s�,F*�����{,dB�����o�=��_,�B�������*����.�U���eL	j) <�n\S��e�b�E��G޺�0��x[K���CG<�w���������W+N:��xa�V����.�BJ8*$E]J�����x$�^���#Z8>
�(tCD1�r����%�&%E̽M%��P�6���
�����VHj,%:Q��J|q�GSi��?���jKt���el�H7�`�{/[��?��?�g����~��߽�_?;��T�����˷'[�dbЩ��j�	��LLe�'��)&�z�h�Dr��5�����)�9L�xxa���'^W��ؿ�f��F�Χ�5�����ب�=��S�s�i��q�����ZX5�5DiKs��F�E���U�|�W�n�(�s^�������>��p��܍��L�3�҇z���r���1�})
D� ̻�cҲ�FB#F���g�T�����"��p���#<�J�[����2�$�
u���CY�r�J�������dm�߱@;}���>8g!l��6������p.)�^�~_�s@	�j����}{�"�Aq�~#�c��)�(rA0��]�a}8��s�Yg��~[.��,�_����}g	ܡ�P��W�@��ZĔ+R�]�FW�.uƶƱ�PZ���:-ORM��S�ҟ�\������ ����贿��~�zvϬ[�;�[�v�(���E�\x�_������y!����3n���������Y)�XNr�Q�ziԓC���'V>�+ioU�m�(�,w~���z֞��K!�G0V�/v��C\K���?��k���J��x�a��^���:�!X���ndyRؾ�I!�祰�/L���J��gG������Gы�Mֺ�N�C��Їrg%�=lјѽd~�}������^DcQ�V
�=�P�M��>����<~�,�>G��Fk�#�2e�{ Bu��2��5����.�����6� 9�S���{^o�y�Oc��^��d��j5�h��"��ui��a`���:�+�f��"~�_�x /�1���+W�H1�>Q�)7�S�� �}ݚ����Ś���G�Ņ�,��x��\��r�0-
Z@����/�rjF�_�=�_�I��2�����A�؁x-z_:N]#]��H����s?���=#&"h,�џA���C��gh|	��חmiAW1"�)�HV�Կރ��G��M7ݔ�85o���}��;�h�^1��8���/~�w>��4�݌R�тz��o~�7�x�aq@h�0=��Y1�~D�O�q���R��)��&�,:Y>�z�]�c*���v�R�2(�B2J&2�e]�-��yJB��Q�C�аV=V˵�-�~~�P���Y�=�s`�{�+^a�y0�:�΅B4�g�������0��̈́��,jfy��q�������*�H�PD4��Aޙ@��}���c�,7VaZh�D�x�Ɍ�Y���&|}�T塘�5���C��3�<���og��G.���?��ˢ����'Ƈo�T�鞙����Wq�vu��1֎�&U��\<�rɬ�v��L�<=l��ΏG��~���&�b�b5�����6����{�"�_�I�&��5���-=����
���h��G<��o�鷃�Z������J$��B4�Z0u���4v���Tϓ.BZ=��b�ڎ?�/�k�,�d���l�"_F�����4ߢ�A{�0٩*Zp�O�Hظ�{|����[��S�q���?�㣟�������%Qyv�϶�?O� �#7��S��DO���\T�|�Ᏺ��p��h��Q���G��w�����xp��U�+�h�vw��C��Z-�,�Ks�RZ�aÆ���^��D��v*�k%���TW0^��r�|}��DI���¥~(~y���=%c=ݶ����B.�7n���v�/Nd%�Y���Z.��̍����0v ��xF_��+dO��Yq�Iy�B4iq��i�>�����@Ź,c�'�=/�S]��ո@��q���.�<��ȌS���_���~������V�`�EG�B��ʯ��OZjB�
�sd��z���'�����)��p���|�q�-#):�����̙��W��e�~����c��c)'=IG)�UX����k�w*)���&�Ox*<!�89!!W`�$�O')�<�W�zo�����!�c�9��9�~�Y�
�(ɫs�sy ���/��/_~�G?��w�m���<^��ZT��4 ���X��.��ҷ$õ?�;{�"����:�dF�g-zr�XK}�L�^cYqx�'�����1���Nr�_����h�X1�1�O,�����/|w��[��T���_�����߿��7\s��M�o�T��RXr�YU��M$}֊����2�a�714�O<?�(������q=��������o�г���Uc���]PH�k��{�`m�+$,W�IAR�bŊ�ɷ��,h%=�7�=ďC�p������V�C笐�^�|��7��y�I'���&��骫�z�%�\�!n�q���1d^h�����},_�(�䓻S�D����g��[^��x����/�QP`-�B�y0����P�ђ|���{sl�og��G����7��w�m��6�n:;��]
�zqmo����+�O) ?�䎓��i�mb,��b�԰�jõQ
�Oબ�q��5�dg�GY�x�_�����G�R��0~/#������>��Ǉzd�J���RH�ڄ��zƆ���?��?�Qu�x��Op���;��7\{������x^�c���șI�
e�=���O����ւVTƾ���-��Iw�������]-J��9}�y{���j���6Z��L�D�B���*����y�����[�����~�����-oy�O��M��^T��R����
�Qp�V���sl�뮻.�p��H{����I��W��"���o�#��څ�כ����x�O4���81���>�+���L��^#����Tq��vi��9�3�_y啗���kg<����4+U��\A�+��зU<�����pǈ�{�ޒ�I�W3Δ��h�f�;�!��� FyGq����֊�W\������n˾g��G�K�ȥ��M���OƋ��Ύ��!�Rф:T���PK�\&Kd�kr0@�!x���p�
	��Ysf��j��;n��N�O�&Չ�+tuu�[�[���w�p�	<�y��{��8P�[a�}��YR��r���a���	����7��E[s,�{���/������*q��׻��X�2�a�l�h;��*�v����z��oG����9.���줮'��kL����d��'-��������u�kf �)m�ɛ_��W\q�;���/���G~�O��d~��#'d)7��<���x|AS�2�
u�}&.5��"��Xg���)/�XY'��/���:�c�)~N��؞����}r\q�f��tW�^+�-Z��YO|wQj�$�?��u�\s�����q^����W�σ�+���(K��m(�������#$R����d��z��>
�f������M�q�^�]y�Ag���l+'�w�����y�{����\saT!�tw/����Cx�f�{{����ng�q�s�����y��Y�U1�r#�6�Y4;�fʩ�ҁ%�v�����+_�J�c���8;�.��{�0fY��9�����<�Fֲ���!ت��n�������:{������+�,����#������^�|���H!-e$��x�\&���*e�|R�I����h�<�`���8a�G��w����}n��n+�:��������ݯy�k�sϽ��q(ύ7�8��;Z�'���|��P��^\����M����m�������ۗ/����u�Y���ٽ��.�&�&s��=��me��]<��O?�l�n���mrmN?��M�������O��O�|����&"i�p���P:R���h㦈������1�&������=��1������ӎ���ۿ���+���}�����?+ޭ�{�����7���#������{��7g�x�:';��	�T��	���|�é%�QU�B�H�5I��3�C#�+_��׿+Z�+C��z��Z�kD����+��s)�����a!FY�8�c��ړa,�����>���;����x��ZI��"���7�a��o=����-�&W4�8&<�x�6Ɨ���g�]��O������{����	�w[�� o{���>���~��{�%��y�Q����dxy\v���0]���WI$CV~R*���L.8����YSa��JI�aҷysR��`F��,,g�rV
S.�=���R*ل��;R�YRuk�4�`pB��RP��;E%b�����y�m���@���x�?�;g�G�F�#��wߓO<��/�.]J�w��Y�f͉(�6'������q(��bի�#Wz���z��Fp�Xyka��%�F����x��h�sSk���^o�F�go����9ȧz�Wuu^�ˮq��R�G�X;���@�}��J�8G������m'ʽUʕ�;*b���Qf����8�x惵�����rg�(���R�RI�zŗꎇ�}����'�\J[ܛ�{T����j_<��{�������C:�8����7��(m�������W]uUwTB��гf͚Yq0΍�DԡS8�y\��%j%dcJ�n��f+��w������7�3N�2Ǥ��5Ǥ��/����&�4��1��uR��'������~v,���qL|���K�������x�~W�Egէ>���ƒ�x≏���?�hT������R��n^�#�e�m��3>*<w�7�d��g�W��H���Low<^����.���,����w	r]�d�Prz�K��^Jo���&��4����@��@�����uB3�;�Z�T��{���;z�I��ܶ�1�W�XfPƱ�~�u����gOs�1�V.��~z�;����y��ٳg/�ے���.u-;^�A5~n��{:���������k6��㸩e�|>_�h��yvM�l��`���K�=*�����54��M�D�%��&��9r<�cw .��K�,�׭wٲek�9���7�%m�?9�l˶�
m��r�i�Q�{O�d�&�(o*������k��Z�%�z׻n�nm٩����ҖqH�M�J�������[�Җ��@i+����-m���V�miK[�2����Җ��eJ[���-mi����oK[�Җ(m�ߖ���-3P�ʿ-miK[f����^��2�R    IEND�B`�PK   �{�Xǐ]zd� K� /   images/0ceeee3a-ea03-4589-bdea-2202a7c6e233.png<zUT\���n����6xp'�C� �� 	'��4hpw�����ǽ���sN��N����]�j�WW���I�	  p�e4  �������u��Bp��$���< h
2��^&'�h�����*kE�g3"��n2'�5�k���}��z��k��Qr*��zQ�E���P�AU.%}�����	�;ޓ�k�EA�������5��Y����� w�+H�UhQ`�����	�dC��_'$�Hn���o�)B�х���Զ!b�`�[�������߰5��:�r�v��khL �t/�����v��K_-)��i7�8yol&�ө�������;�FF;����d�^#��D�a��|�����i�2���O,i�B�K)����SJ���	�d�`�-ǺU.��I���_�a+^��G�+�X�Ǹ��K/R>2��W8G��R�%�.��*ou�G��/�H�9u��{<i��'�G���'�*KR���k��n3V �6\�;l̊�n��K��x9���r���9�/�J�h�~В,y�t��J����L��H"ˊ��r�k\�}ff�ƟgVH�a�
�q�,T�l_V]z��)���<�#=�B�6f�z!�]&�5��.;ޤ��V�������r�{�n���������)Y�km��~��$�� �gz�����̸YN�#�f��x��~z:ٞs�t4hӨC|rS�ǅ�9?�UFr��?M�?����|�>\�5En�$GF]��O�=�_-;���>|֧=�!�����X�38x߹�s����SǮlћ���ۂW"K��� �r)��pﺐ�9��_��vw���ֶ�NW�Η��G�ZVe��?����Qۅu��|E�켙Qz����̮�+N{�%��U�ݪ͚D��L���Z"k��Ǆ�J��%�k���< �z1�*���Jy��DͶ|Z��1��3��
�ٴ�d7��[�7�s��y�j�sL�kH�\�o���H8��t:�5<�+#��6?̮>`�H��&)ο�P111�WwN��ڧ���*$0&}h���:%��d��d��۱�5���a쳨*����'�A!�+��G3�)�t��]E�0G�4|�@�����]�=�'n
3ާ�����0c�oi�-3g_����Y��8;q�t������Bt1pVc9#⣙�tӷu��p&��������(w6>�T��i�
��i�|4��@k�lHش?m�J���敒9DX�\N�(�
<B��T0�+k�.e���3��	��!���*���l������Fυ���w�o�Yz�]O���)3��P� �������Y�E��a�k���VUq��in(��L1q=�5��s��,'{1��L~ ��d���<m�t��n#���y5��ξȸe�N<�B�x�h���0M�}��]�C����4�|�ʯ�;~�\���<"1F��0���(����cCgK���;cqC�d�����5IZ�ln���_�Q�����Wnr����Y"�ٞ=�%���������g�)~-�����O���%ȈA�����cRdR�}t � bn�����8U����d��>��i�����IN�_?!�}Â)�ӃfN�j��z��{	�E/�vj�-��gBrh���F��FX��AꜾ��h���G��I[�l�Dds��if+�Ṳ�q��>�l^kE/ݧe��>��߀e����·\\�������<�!���GPeG']4��k����F����?TE-ݐ<8'k+s�0��Ш�����x]j��U`C����]�D������/��M�'��⚊�y��26\U���~@
ش�+K�S��CZ[w��`n\���p�A�u��h�x��fcƷ��_�c��N��!/���*~G���Le�Aċ��
2����!"�0m�Oq�ّ��o�v��'���=�r�1Fحt�i��BC���يO��]sB����n��@����1��VМ��K(�}������	�}�(��V���%t�p��UI'�^�P�7-��K}�:>bk������Z�S�W��T��sW9}���}#�>�~�����Q�bР���bBt�rF��Z%~2�c�����������B�!
ؙ��μ��pu�S��Ɏ�PF��Yۅ=�5�[�e�J�$����sC�(�"�tc��2'v����%�A$d�9�z�����w�TmE��꽍#�)LP-��>#��W�.vw6=D���
	~ �l��"�n=w����p���Q��Q,��j��LK�7�vU�6ϔKX����{�����3fݥ�VH�����W�+�s�ȵ_G���fz�+L7�e�8�n.�Ґ5�2���#Λ�N&-�Y�P8�CC�g��|-:_,��{���4�zb�Ð���Qң��P���I xP��� �@��pR�=�� �Pm�3��|��l�Qd��5чV���A0�}�v�{wS�� ��jX �)�s�e��"E�"�����kF��/Oi{ �n�*$�<氿>�O��4Hg_!1�fc�U�8�c��ke�R�9)y�(�6N��T0�tUi�ܜv��]�e5씪�ٓ�f��%��,�b���Ǝ��/CJ����zd�(���!=����*$�G�kq߄;����s�r� �QZ�V��]��zE-s9��8���ɛi��侮��չ'~�A�s3�TU�����#�(�G)�-�K�=�m	�S��S5u����U�ܮ��T�}[n{���H-�Yc���~�ը��{�����=����\�����3B-����RNB��_i�J���8v;*k��g�ܶ[����AU;F�$]���2��.dA`�� s�w��8h���~��x�~?Z@�뚸��\.�pD��O�����h`���@��X�~J��K����|O�_�᩻&i�1d��>[�7�:�1�6]�bW�RC�E|6"4|���l�tn�#]��u��J���o������a5��/����o�{���-i�{nu]W�; �z<	���_��(�֫���F��nM��d0��۵�@ ����ˁ�2�v�t�Oܦ|k)>��+4� ��=��o�/�%��~���[�92��/]/{N�ק��}���ވ�&���jwP
��dm(�AN���z8����%�Q�Aܕ�����@�/�U�s��D���gK��N�����WL�G��un���!���O�U��f6�2�*�?`�
ui����^�q�*_���ٷ� n1M�	O�����Y�|^[��~�R���_1�~��~��|�;��bP���"�g��訬��b3,{tt��� �O^)1aw���rнvZ�q� Jʗ�)�5�+0�n��y�4$�5���Ga`�Y���H
e�5F����~<��Z����s[�a?����̴�P�^{���>�r4�]��f�+�l��1�tߖ��o�W�{q�����0�Eد�?�$E����.��;w5�R,8'T	�?qepF��zf�!�UX.�i]Ͷ��S�/N��{i�����Ǎ�����sEc�7Za	����B�	O͐�Ւ����=<J����fE���s*�U���2�
�'�N0���ߝ���m���A��՝~���~���ߢ~M��ņi��j��LŊ�k��x���f��{�s|s��Κ&�K�-z�$/�g~���T�5~*�+�gr	����>a�܉b�*��M�J=�Ӊ~��^�7)z�f_��$�����5������o)�Fp�MQ��N�B���u/<��ڬ:z���='��?���J&�:��8����U%���� Oc1c]�O�z�h�/��LŶ7�h�\!�~�7)�II����"�����S����y�J�M�`���]�m�MN{�xh���Z�s��ƚ�u�������/�D�r��s�2�`S�s�7c�>�	ճ�'�}S����Ӥ$�����J���WLV�����5��t�����K���x����q�kd8U��4�?��?�O��¦�T��_�L�:�,W�^��l��H`T�3��P7d���3�����(��"����N(^��S�Q���+�K��������⼋�Ѓ%��	�y�9����݉���~�}oܴ�&k�;\$rw�J�`S�����A�ۯ'�u��n�|^ú巏�㧳n�k`�'��S6fV�x�M��� �����v0�ړ���*"�9��
ٸ_��`n���9x~ �e������\o��:���7�%&^���k�?�,܉V/�B~���Ia�3�q�=N ��t���=������-�dU�w�$c%���>~���O����c�)�#�O��4���w^�H�R��I�Jq7�@a�E*o��u"�E�F�L����̬m���M~���;��J���S0HiJ�2���lB���b�����OW�Lfz�g��T�m��ԏ��	������-����;��Ґ�(H�I`�.[�%���(�<Pr��8F�"01��>�/T�PCS�:�b���(x��[?��I�������_��5O�)����� �=�m7��H�y���c!#�Xm�p�P7<`��EPD�����Cm�?!���[1�.��^���l����p�6� px:v�ⱡ'8T�,���r	��X?b�@��@��&:�̛�L�*�׹��4�J�e$=�{�
:~|g����|�!������:N��$a+�9������*Z����j[
Kg�����}Eze�j�lM������B�Ϝ*�I�@=��6�/�N���D�W5m�}0�� {a���W�q=?eHP`9�!�����VQ�?����*rJ9�q`O,��L�H�����������K�ݱER�a��@r�ȴy��P^H��`P_��u�������I�U��bD@?.��^�Mv�wN��n�p���[��a,� ���B]X5���?�qzP����I���m�wcK�lE��5���OYh�,e:+���靏b�HA�^eo���ybW5X�9��YBޑ��T�Sb��{ni��z�p_
R�o�4pc����i�Z,����`v�d
ėbv�W�!�4�wj�N�*���y���3�A���[�/��&���fX�d�oC4�
���+2Z�B��$R���
 YSu��P��G��L�m�*�+���mVp�]V�ix��%`�/�]E�-"�w��M��< V�7�ȣYL��k0�P�g#��ڌ������`~o4�c�0q#Y.�4z�������e��� $4����㪙��f��zǕF�S6E�)�+T"?�Sq�P�ߚ�(��l�j�����{��w_W  ����K�ru���-!fjm��18��="K����ڿ���Q������k�uFDgD���?j�KmTk$J��	α �X�����$5�1,7��~�����d��]k�����)p�\�n��.������F�{�jƎF�d̴���mX�dvg8�����3WHC__!�ԫ�[��[�	B+>E�2��@��3h��5���'��f�}J���zF���6>/M�9�ϝ��^M��b����[�j9��9-��*����Uʥ�+M�J�m�l�U���&��7�䢺����P�b&�.��_�1�N�y�>\�z�9.[	���ǫ�K�<�����Im��:�m��?�+#'?Q���ǟ� �J��OXgv�>���{9��=/q%l��C�f�:n9�*)&]��'�j�LNz!Xkd�&me�<Ԉa�J���O'��O@��4h�wL���ZYխ��xQ�C3�.#QT��R���ٚ\3	\Ԥ���ے(�����_�h�
��}c���U��]�_���Zj~�jr2eec+��d�B�:B���I��^�$I�#� �N��0�fe�q��gOT�U6���� �f��]ۑ���}\���b����:o��ɗ���fb���\�茆�ژ!��Y�x�������P��?8����nch�i"���շP�Άh�'eP{��̻����{8i�wa^�b�qw�vt gls~n�����@�7�JƸգH�_!�����t3�V��Ȏ��T���|������� $ ��r!�8����Y�X��;�7�2W"*���+]�Ի���2������o�P%����C���ҍO���6v��V�)�	����X�$��w�<�l�/�}��h2ǟ����ӛ}�K���	��Ҷ���]�(Wgf������Ѓ�	�zmmu�%T(����F�sY1n�O�+hb$�$Yon�w\2��Y0��r�9������=m��������h$���Ğ+}���ǭk�z�Y��Y�+Ĺ&5P:���H`�%r�|��%�sݛ�t�gw�i㊗��]S�t�B�A�g^M@�'��@T^$�_�l� �x8=�"=M���w�%Z�2�Y/��O۩�'u�:V�2�U8֊���c�v��C[Y���:����0�����Xшo_�������Q��<���Lhܦ$ad�{&���w��E�<��*�!H�u�|�^��M%AH��7gk�8��%{�� �o�̸�)�����	��O�	���	����)���@�����A��A��kD��>�t�m �D��8�A*�m&e�J���<��c��U�I�p'<��]�+�Y.ܤp+����MB��~���=�cN�3�������m\�lkB����W]�ǩ�P`ӼC�gЈVֽ�&���b��p��.�<ߟa�/ۣ�6a� q�L�o�A�L�^t��y~��e���������?B���:��?#;
_NS4{��/)N׫��Sl�f�'M�2�X����<!���ݻ�{�F�W���n�'6՟�����6�̤N��t1h����e�j���^�d�"r`xC=By��K��L|?s�����卟�h�xPuR��r�}��nc�0;Y�m�	!8�A����&���O�ߜ�)x��!2�:������=���7{P-h����bШ�h@41+��	`���}4WF�I��k�!WhS�L���}�9��"v�[��m���Q�6IU�m�gY\CT���ǥ�ĬG�)B�Gs-�D%���єj7������/>a��/�:��uA��
��Y�3`%��Rc_�x�3{��d�Щ�r��p�i�XV,�L�ڨ.�[�n�r0TS���$�'�x�����]�	O��w�\v!�FFDx�^�͂l���|X&N��3���P��^|��؅��:ϑ�\ ������ �Yq���-����q��C�J�z�@�7�+&mk<�e0��~��t!�b.�OY����R�[̘z��p�&}RUm/��ҿh���ߟ��/I��_p3$��#��Z��&'p���ɴz��o�s"�X2�)q��z"O�)�.GP��X)m_+����'G�u*Tŝ�kHҭ��.�mȶ�nX
�gg�P|���,�%:i�.�"����i ���3��qS�W����4�R� �v���esCd�~��w�.��u"�=s��bv�NC�  �s�0e��h��˙g�h�� ���8x*���Ծ	���R׊�5��᭦�{1g�jֿ����_�{�Ǥ'lRc�z�#0-���Q�4�41~��-���)��.��������jFZ}RJuq�L�*`G����Ҫ�Վ���r�J���9�ի�h�������m)b�/u��.�<��6��2�BM��-������s�O���U���~��͙/�dyd-����[�Kq�mXM{Z�/�] 52�"�T��-f�\����J�k�V�k���U ��C88/u�H�Ġ�@��y��n�/��(�Hq�"���ȗY��ea1B�4lOeu�g�kJ����s��͡�8��"�5D�{�����+05�L>M@��Dy�e�l�I
�ȶzw�����A�����a��{o	�=@U'���Sd�^�����ytz_�_����u>̷Iw��mћ��܅
�l9O�sF�����|5�:���	{V豝�A9Z]Pg�{��~�C�Ƴ*������1����3!��(>��S<WcQ+q��c�վ.Cy�qP4.�x��ǈeh^qU��w��Ƀ�a�rN�d\�%�3�D��]��	� �4��fv��E�c��6�^1E��v�	��_�
�@���r��l~��h��{�Ag RP�~'�r��p���1*�W-�/
�(<Ȅ�ʐ~�Bu�켓� ��hx'S��A��6;F�q6�E��>տ�fUZd?z� ���H�E�9,�GE��S��$]/�Wd]z�{��¹��Ju�1�|�9>���U#��E�����?��R!v��%�
ٜ
�hE�"n�漱����5T�-�ٖم�ݮ,)J�ܨ:n��$�A����h������vK��z�GS��+&�J)������z�H�T-�Dج�4��3�LN9�u��`�y�
�>^P<�I&7��/��%:��F#���oɒ#N氎��d�۹Zs>o&�4�#�'A���)�f�*���#<�Ͷ�m�w����?d[���8��ƻ�U�ET��L6�J�D�:go����&��[����(�� �D�E����7�y�P��;�Ks��kn�m�*��r[Q�Q�"dH� ՙ��t�_2*(�:��z�n���B�Qi�N-�;B}�ژ� l0ZVnD)���
ǐ�2����[�;[�E�E�,D�Õr��,�%ܸUx%��&�H��:�e굉������'#�X<�7B2�����R����K�Xoo��&,�T�1(s�<�hM������+W!R�g.:�O���";#o�~ˎ���a<\�{�iP��ś��<3;�:�=��nzg8l�aC8%Z�*�ŠÂ���o�����4�&�·��X�*�㢶B����츉�˧��lo�a:�3 ����T�;�)w��C������R������y���Wg����.�n�&<�u�^���rr���zȕk�8�|S���/�� <�w�L�Y�;ӛZL�)D���k�V�����\������]�I��ӹ0a�t(��\�j!̾��\�x�?�G�i1d�T+(K�<I�,�i��w}���k&G&���P%�D�Z	��5˘�����g4c�<�۔c�;0)S&�K�;�����<���Q��ϻ��ZTt�]j��J���l�}|��\��UC�y�Z[�Kժ!�E�Xhucw4%\2#"Al|��ƀժ�.{���q�L�/E.TC�oI�Z�x�b:UQ�1�!�)�5����DšR�*��_�z��$[�)���M��1n������cbP��4��
h�����V��"ǜ�?}Ǜ���߷ߨb���Ԇ)#���j/�����ٹ.��>�����t����Ƌ���M��V$k։�$[8�#�7YYX�z��q�n��L��Ɵ��.�?��>B���s�8l\ϧX���ZBb�$�]�8T�nLm��'|~?�ʝ�K�����-��������u[�X�6�Y����[��K�m�$)��Ȧ[�'��c��cɬ8f�7A�W^�|��p����?"�WՈ[I�$�2�w3s��a.Xl�u���CPl鍍�[���͂Lf�����Px�Z�������;�4<q(m�o����+��%�w����:T��=�9J�4�[v���@M���Z�<+��#	�Y�\gzj���;��%W�7���v���Z�����gaG
&��o������uo��\�*�Ci�Sd�齅�X�K�x]~�k[Ä�������pa8��'���;����J]`�}pF�$k�aӿ�]�b&j��ZHJ����[�Nj[��{u{����m�s���N�Y��&ݙ��qw���x�2�Ѭ)��W���g1`KzI�-nzX���_N���-�#�?7j`��r�/[�D���\>�u��L�Z�13�o�B�9.���h�4�$i2Y���"�����,C�؉Υ�-"� ����u��p���ꢁ���g@�������۱�`�=I;���&j"����NmJ��am٢�2WP�&gr��#�2�D<j H�(W���B=]��?���Nf����/N;t�"���t�}�tOF`��S�+jRԸ���d��G�����i�H$= %Z�}u{c	M�0];RJzD�<S���u�v�Q~)gʎ`B$��Hf!��+Ֆ^���̠���_=��8ABL���Bq��zb���R�W�rImK��� �WpK �=��c��I$��3��	�Q��_���z5ʥ�4辉@�:,J��'&bY�A`�xr�s��sm�hD�&�+9�O����tk����q����Wr��`~��� X`������֛KS��������������)��ő�x/eV�C+,v� ���*S��yW��<~ �4� ?�$�i�C���V��w��`�����Ub�`������Y�%��}	H6��P����B,"�G6��xW�C����'x�H�T�����e��W�<7T�GN�����'[�caE~Ks�3�JGN��t9���3M�_Ռ�-�y�;o�S�������zC�c"k�%���6� �b�e��x\#�� �q�|��9�s�]��eM�fV�E�/��ą?&s��:U%0Q	e���F'�ڇ��U';�C:+��wބyMy����*Y��|ǫU{L�e�,�9e&�n��«4h�&�4Rݴ��&�K�N.�%�Z2����\،�z4G����lk/V�E��e�s;�
U�����du�`g�sҾ�$�9	\�������beJ�P;ߣ�aml�P�y[�#��������_�a� ��ƶ�s���� ���n�
��	���nҠYD�OY�aM����y���u���>��f<ݽ	N��Y�&�����eq���{���9O����(���&~M�� �Ѓ!��?����*��!Ѷ#��!Q����V�C,H6�7���0]���ϭh�h�c��9���{N����?�����h� �z:57Bb�Dy�D_%�8HB���Ys���ęS[JsY���@A��O�^&�9�+�k���e��(�n߹De!*���-�a��58��:�C�~��p�fiF�1�1�1Cn�������DJ�m!лTWN'�,����8�>���A�
1����c��񥧧��f2����e��I��������"���=��!�� H���=c����rj��,����|6m۰�8!\˱��Zo$�;G9����mmy�cm�^�QgHTxIƕ���N�8	����˭�Uܐ=�N�>le>�|�i�̀�ާtt�x�7�u�<�o�es���"C5>��h�c1"Vo�l|M*��q��wk`Q /-���$�y�w1�@�����Y+��]w/+�� ,��s�׺5)�}5~T�a��i�o��hH����?�b6;���OL��5�|C�i7X�<��Ϩ��<���+?7�kao�`D�)@Խ�ː��l�?׿��G��_֎�A�PAD��Hj�#-��-�xi��3 �'�H�H�Y�-�"b6�y9@��=��zW�A[O����P{f�)���*¯h����3�B٦_)�4/�E2m	?�M2�h�#d♍�L3�����G�7㏕2P~.�3N	E����������ܝ�B�y����yO�TA��z�/&���BP�d���u�;`v_7]|B�I�]8��Xn�2h�87�{݀�%�]#��;�����ʈ�0bA�� ����#i�a���D}?Gћ*ɻ>q4_j��^q!��?n8x;WR�@!o��(��B�Z��hh���_�|��§r�/Y�(\���i|���S#M��5��O#m�@} 
ܠ���E5�������'x��\���'�y��̅y�Ɠ�ѧ��d�>��*���&�Q��tI�_1���3�`;������B(�:Y�P��`�<[�NŘ#Ή(��op��Ѥ�y��M�M%�j�w�Xۘ7֬`����R,���/Uk��0z��?���wD�0�V�~i>�"���/W�S[�?V�DHBzs!��5�(v����\������fDh�PG �������xۙ�����
�WR�+�j ����x�Tt��p/�$���������ĉ��;	j���j �⎸���ƊweI����	��k�X�13�\��ݓ}�
�_w_�����=���HO��m�v-�S�-�U���8I�N�����Ln�
ɭ�s\d�ɸi��`;`�Y[�Gji��ґ5�*��o�!�C��)�������p��a�z�Jز^%ʔ� �� �.��;�X�I�Q`�G
�y*�xf�3B��C��@���%"�<>ܜ���7��MƮ��b]���o�m₌O�<�A�@�g�Z.�u1z�����D�΍�u�S�fo2-���I^�R��t��0��M����8����H��h�ff�8��<�M���"v��Tؠ���f�����z�՘C��Dٟ�xɡ�oe�����paRD��W��1m�����* �k��<�.� �wo��.+03�W���[���bUQ�g��,����T����џ��l�-�+P�	�x�Ar1ЀBc��1���ˏ�wJ�� p�oN9+:@���8��RKbBN7�N+ӿ�crrO��[�=.�w��d(/fj�lV��&X�;�ϱ��ຉ±��@�;�D3Y�bCY�L�)��@Pa��6*�S��[d=#�["���R74�����&�֦$I��1S�d��[7�;t�]t�^��7B ����q��u�N0,KS�\�X�(�8��C�q14�*!�B�^Ϧ�������ę^I�~\,ߦ�Sǀ |,l���[��!��z��[ɲ��JS2��Ԩ���L�x�����6>	;�cYX�S,od�HK�0�i��ᓎ���o�m�Z/�ӻO-f�U�F�c�7m�����	����;YXj�̓(�$���H17���x�ӻG�.��Y_y�vv�	�tww���mrTRFq�+ι��nY�tj�?Ŗ���uY�{砑y�o��6�1��"��5�7#��1Yʴ�	��ϙL�x��+Q��&+��Z���Y�=�3�֖q�K]�*:I�����$!���t�Z(q�oXI�jdB]t�0 "ÛKΊQ߅��	jɐ�>�!Tz���}b�d)�`3�]��m�Łs\��=��=��e��m슧ў�  ��vM��*�Jҧ���'C�y\F��F�*?r9;�uM��I -v��R?Zy�">�IY�s�ʍR�=�-A�<�?ݓ���)�P��vX����{��1x̤j��Z�c&��O��{�j ��c>�4wp����Db�w]~��"�;j4�^��r7W���t:�0@����;y�o�/�xzX«��J�3b�v?�
��Q�^n���8��8  �y作���5H�TT��\U��XNym�3�����k~��ƏwC��J�H�Ny����|�l᪑)�=����'V������ ��^7cI�ǧ#[e��̜�O���!98p� ���欕�`eF��E�Y��z���b7�(�)���1Ż������ԥ�~4�� ��$21{P�[��_=��V_8�������%����#
����b�����3?��.�Ow@�^���H��t�޶��/L
dW���_��I�:��J�.pG�}��`�eQ~3>�/��A���:Y9��a��5q�Lpr��;&U�a�6*����.����a.C	��u�ջ"$3"0�2F Y(.R�^*��;��+�E�h�|��7϶��]-��\y5Iư,O��2F5���"oڶ����P�/����=Ah>�j%��9��
ճ�����T�����C1�31�w����L!�����
l�ɚ&��s��c����R��D�<RS��:�wc������W}�Z�ꊲ�ȁ��>���T���1_�~�w�Db��޹A�v!<TA�,^<E��BF�>ZX5�k�~Cd�Y$�
wÎs
f��&��@v���v��s�� �:�+�Β��,��yw�5�xr��G�a*+.�pZ:�B��/�?"��Ⱥ�F�ۋI�,���xs(�0_J�v��;W�3w�-Y��\����������Opr�Ao����5�čM+�ѯ׵�P�^�i|�puc��VϪ� gd���������-�9��ɗU��0|Co+�b�o�2Avn��ʱ�H�$p���5�w?Ұ�����+�
%3�B�q\i�>�8�@��ꒈ�q��G�N�sYA��5�(�"�Hy��l��Dc������9�b����>b&fT��Ȧ2�C �(��g�	�
%�$�襒��QU��Sد
���K[�a���p(2�gr1 (��z�=�9�Ш��&�H��D1�������-��(�".�ءF�� ˋ�و��S�W�P��������m��N����<u��Wu�x����H��S8D�܏�q�;f6�4�v��հ�uA��%�4%5H"���= y�1���������*����Eo\���uә����I�F4�"�#b�k���,��g�f6?�;U}�j{-�W�� /	�x�P�nĠ�
��n'�+���\J��OQ���q$"��$�S�J�8ƳD���C�. ~�o��$8F#��/r>󞆫�ſ�A��>E�~K�;���&����Q�ꛡ?hq_�~&s$�V��Y�|Q%u�i�B��hM0ۆ��"/Ɛ�O�'=��Եa�I����J�������e��%�ҀH���EM��,/S�?�D���O'�AO��g�h˔4�A�\����Y�b�:'͎����'Lc~�3^�D���G_�����$�v�OC��-�����?���@]"��J��<��A�����q�Ue)s	p�HbԽ��w>Wćf�/�u`�JA[w�o��u�����4�%�#�4�.�RJg�-\/��g�Q��{�|�gTN��[�)�
�MҫA�9	���c�W�zӎڽq'�E;HG01���-���+p{
6$����Wo�:��MF���fv��f�4»Őh!�s�g�A�p�IL���c-u�N�����)X'k�ȖYQ�N����7������7��B���R0z��	�:�8F�o���ԕ�)��keO��ӱ�MV�S>po�/M�J��mJ	(U�ӎi�V�A P�N_i{ �H!A����s�;ć_t<!��ƥJ�3��_.�$����E��:����s>�S��<��+��)�/Ma��{qX�1���e���ڧ��G���.S�>&j"��~[�´L��onYu�n˺SG�0����jG_����+��#����ی��N��t�9����X����k���g�ĳU�we,�ڥ��tM�ӾV�{;+ks`�h�K	?��[�U"u��#| z>6m�}��z�]������)��ltĉ�O��I+t\ac&_W���4��-U/cO�pܜ��U���J��ݸog#=��s�Bh-�(�TyuyS�@��{����BES�l0�9OBPqO�B?���5Kh�n�3��B��Ry���ѴX	�
/���w�VB��"��SY�e���t�8'�UG�I��W
ζ��H������#v%3*�k}n�coO�j�g�*ptTN��"n,�W4_��;bª80������[�D\�$�:��Q0����S w"i�x������]������X�-um �}Ko�P�b7�~�3QY6U���P�z��R����<�U� �)\/K��w�L[}1A��9JM����y����=3������_,�[�#�w�Lm��H�wEiV�8W^	;�2�ն�GN臚f��a�>��(چ	�������'���r��~��I?++����<K>j���O�B}iW&�ڶo)$�|�4�۩�;Š)dc�!�j}�vs����W�U2�=܋$ooL��4��+TΡ,݇eC���|Į�:k�5�I�?���Q��o�� ��ٯi�������g�u�&��՝���cL4���{ն��.n��Z�P�䉨�$�P��vzK�r�D�%��U�f�=�Ps�~0H�?�ԙY�����Ȝ>��#|nh3u)�'u\ד3lr̽��g�n�Z~k� �mrXWtߤg�0�xH�z�w;�7)�+ pIJ��: �e�ypG��޽OI׫�H�\(�'���Ua�S9L����] ��J�o@��
]'��ꊆ��Ǐ�b-D9��~�)
쯝!�D�XM�o�����`o� �b_K�_��=�������NQ/�ڰ��ķ�T*�WS�0�s� |@���Q��T�kTJ�$Tcq�?�����=����S9�Z]�[Ə�����?q�.�%����?�Dwǎ�裏&#�p�F�(_Ck֖R�����9ulv>?��Dh�J*�ї��VBy��>8k��2�N�|���5sf�|���>ӊ�U�.�� >f�u�LW^y9u�O3N��2�F| �"5�a�z��gì7H55u��2������?�T���/���������C�a��.����A��.a�ʕ�F�U����w�Ü�
t�Q���ߓ���./��t�J���~��ʶ�;s?�0d�զA���=���1*�#�1�
�����i(p����������ߗ�)e��c��~�q*-]Cy>����0��Ր�)�z�L�8�y�B���T�R��ǐ��<p5)�*���i��/����P߾}��4z��_��W<�x���P���V]�VZ�t%�0 w�o}M	D3��`fa��ul�[_���<�\�p�$����@�^�CѰJ#��B��Q��������~���|�̥р�}��%ũ���f�z��<��^�֮[Eu5���ϟO�7m���uDF-/�D�FO��/���n]����x�*����Abp|>8v�}�������$(���|p�Y����}��E�6��үi�UL[yL/��w�U�6��y�Q$lq�#p��}z�,Rn����䂿��Rԃ/�U�v��m�/嬟�d-� 6e%b��E�ԱS<�
��x+u�`�r��d�9_�IlH���?�<��xz	�q�i�����oyQ@>T��.@\ȁ	��W]u;s�>7��i�TX؅/YĻ$�#%+��d�jJZ^ڶ��:u)�+����� m޴�����iM��j��ch�"|��5k֌��%%	�*/���ϙ	����M�\{���*]J��EG~F�֮-�Ꚑ]l9@U�:*[W�Lⴶ���4�P�+;Ā���9�1 ��G ���'��'�� �����6��;Z��m��+)T���nZK�C����p�x�h��-4w�����A�!CQ�>�U������j���z���?����W��Fz�����30(���ѣa�E�xS80�z|A2<�o��CǮ�.�3y��(�08�4=L��,�mٲ�����8�^�o�2oPC���1�%�/�0��0 ��\D��y�ƏF�:���ҕ|m���(&-_��j됴.E��A���N��������իv�m]�w N��JQ����W��9�|n޴�^{�E:��)�>Y�a-{ư!(�e�__���	�-���#���C�zı���]���.��
P���JgMǃ���Ac�r�F�֮YF��WR,VE>R�&ȃt��o�<o���~D�5	��۱�0�#0aT4���j�.��K=�#����?�����G���V��+nG��䥗�kdz�s�"�t�T[g�דφU[Q��8�$�[n���)�{��٠[YY�.\��Q�F��(���о�m]t�>˖|I��7?[�N�hU�reo���D�)Z���o;ڴ1D	�K7�p+���y�>���|��t�L?�}l�#p�WΙ9�QW�Ϡ}�G�z�^}�?�����)�{��tđ�r����5�LD�A�QUU-���@���ʫh�I� h�>�(h�6<�r�<��s,y�a��T�38��sU,AL��+3n A^���i$��IR<
�~,~���h���޼�i{e�?����O�K��u�_�=�Ye.@q�Yԛ�C���#x�k��o��ϋ��a;�@:��Q�1��ø��&�
GԾ}7�2�H�D=���6�����2k�!ھ}���;��4v�g�}�����w� u�������|����u�d]s�5�[زq=�{�%<�7u+�H�W,���6;�;*�%h�7�(�C�_������^�3N��y�OӺ5k�8�����r��!�Z?�Pv.��%]L�J����?��:��R�n;U�l�bҜ���i�hݺ
*��Fյ�}ޅ����{���w����d�>x�W^y��}��!0����@rA��u����LI�C��6�	~�@�$D�'�Q�C�(C�> ���K��oSUu��� !=:\���7�J$��������i�?�۴v��'N؟ƌ:H��'b�1�<�����d�Cy��dz�9:���q��H��g猷�z+��C�5ft������4�#���nc��*�B���4�d"BK����D-�UUo�H���>�c	2� ���Bk�ld�m�Y���I��'�y��ѳ�=G���6� ��Fh�$ZG��O��舩G�9g�I5U���I2'�u�z�Ek(/_��HY^
��Q����P^�*9�l�!�4�����p}��]v�et�����T^^��@;�� " ��. �C܋#�2�[층C��WD
zUvB����:� =OЖ���ʸ�����S�~�bfgVt�_�>�Y�q��i��8��<�ݾ��:w�gy�5T1o@����H$T1x�l�k�Oe��y�*� �:�;�<*�ѝz�!��1���#/8}`�=��C.L��O<��:�(���5�T^V��!�����C��C�E/-Y���7�8�|ew�i���胏?�pK��>�x�6��7��ɼQ<�d�w��t�Yg�AÆP,RK�U[��r��8"Q+�d�^Г0�F��H�G�������/���x 9^��	��#!�����R��X���D����M�雯>���j
�}*7�O���─px|D^?8��L���c��/W�w�t_��8`��7�?%���[����U�D�Y!Ês�GdL�rN/x���ٷ� α��T��OU�CN}�ʉ9��g_PM5损~��0�í;|�P'��|0���do���v��`��F�j�����G��W�i�F�rĀM6�~��!�P��9�D����#�������z�x���4���l�>`�lauG�M�<�N;�T�ٳ;��VQ2���3G������CAC8�î۷��	�@�g�[(��u xб#�� T]�u��JE/|�����2�2В�g���i���H�8}-��y��L��iS����T����={��h���>�d�@8)�'ڎ�$H�I�'6��Y�(��2qm��R�Cg$�|�53i�hX�6�PR{�N���R�G���<<�˚�W�ʕ��r]�̰XK��
l�f<�D�Ka�+m�}%�0�2&^)�g��� ��&��NU��ţ!WOD� n��#*�ߏ$��j:��{��, &g�M ��eRׂB:��cXY�=��Gh^)hc�n������!�O;�:u*u�܁�-�џ��L��s���^�U�V����`�׏��Z�1���i᢯�w��[���1��T �G��:��?�A,���S�$vk����*C�eu��WL�,��փ����C��q��m�����x[��o� F�!���oLd�|����|�s޹��c�q�8 �A0 J&����^ �-^�m߾�>s��d\mg�yLQ���@ｿ��a$*A�i���z��co����D{x�n���[��7��&/��A[�L}�	���:�Sg� Ε8e�Ef�.y�)�+I�dao0�C�����p�ް�����"�8O���[{ђ�幄�D�ޭ �,��G�^Y�2�������	��l#3J�F����R; ���<d�a�MR^~'�<�p�/Š(�|\���\1̲8h�w��s�,��j�5���!+�|�|��ǻ�5d�`���0)�>E��	�1�H�_,`�eH�P�����4�7��G��)� �	w�ѣG�ĉӞ8�M�3�H�~�U�Ѕ�ϋ��%D"|=p}��G��(�+��������.��w���3�������z&h��iC�J%��1�DurMP?y�v�F�;�S��Kp��xRe�D\��bٚ�����Y`c����r_�/�#�s�^��8�3W|'Z����8�8Ydd!�׽+�,���@�%ͷ$��;��v�eW�FԂ'�+�"���) �c��[v���󥾄 ��&� iJ�E@[ȿԻ@_�x����kQ�I�O�w�}��_J>3E�D2�>#)�� %y����Qu�h;�б�<� ��GT��~��ڸ��~w�oc+�?��G��]��c��ǜ9s�D��_"��%0����!�"E�eG�>GL�E�@�{,ؒ.�	��
������vR"w�ഖ�6����$��a0 �m�F� gܸ���v���D͐ÿ�b��z+}�����/2^���g��#G�y�����Z��cၫ'4�>"�ҧioJQ�f;��B�(�f?�R���������>��:�*����ۧ��L�j�}t�Z�P�|�  �F.�s�'1r�}��/@+�X��~�i�jc�$x�#�
-����E��sJ2.NyN]C籱�H�~�|J�|�� ��� ���Y}7%�,��]zۤo�|��ޘ빂�|?�To��c���CGR
	�L"V� �RA��ku�\@E�=9
�5}�"N��r���!��&v����O�;�z ����pA�0�y睼c�Dh3�;�v��(�`d�1[�h>X� �ʐ���?\XTpe��i%�������a�hDe~T@Z�dᓉ*�������<0T&����@�2R�"�
�P���q�����s��>���O*߾��"���@����j�"ڼ���*D�f�Fzo�'�d�챐��Ճ���k���K�]c�	}&�4�
`�J&�l�dLu�_^�e�B�H�Ut@����:��6�_�r�����
l��,$2�B�0�E��.� Y�t�^��m���N�Rr�>)D$�+�Q��Y(	}.I���`G����+�0hp�	����G�+���@G�7pu+�G^�H!/��F�n�����;v�	����{��x�ͷ�G�|���#.�����v����(ʉ,��C��O�%d ���� �%��HLͿ�c�\�^�I&\&���ŕ�`�֪��)��,&%2�q����ė��q�G�|��CI�!�i��G�d��8�A2RaZ�v)�Z��k��^Z�v͝�1��*�����5�\ku�d��'ͽ+%� @���g�E ����`ӵ^L^	�G_bl�ѩI�����'=d_
wX�s�w𿠦p}�nF�`<ڀk�}E9�3
 $���e"�c�w�L�_��SG��<�h�����˞���~�/���P�}w����x�V1�Ȅ�X��=���~4��IdQs!Y[�s�X�9p�>���y�F�����@�����[hђ��������@�z!�3(]��t-� n������@d�q�$�t�v?��

��5k��m��9mz��U���f��(���D��\�.����f��Ź�q��`�|�ǵ�L��~�v �>Ĉ�E��^����P���6Њe_S<���@�JK7л�>J�����r�	�plk<��L��"�Z�k�a��h��������ݔ�1������ୁ������v2V� }�<� ��y�E�Ƃ$;H</�{8�%���0�b?��1��)���� &;F�%��*#��L��DD)<��(4rd;O(h3�Aa��]��c��㑘���a�d�v E>�z�J�HE��&��7n�rD���C&<�z�N�(�x�����|ҢD
6b��kp,j���+�p�1��9�}�)]����B�!��E��cA�� :�J�CY�kd�(��nW��1.���"�4�6��5|ݧq��G��k�2x�Q�V_���߲ʋ�&a��	m� �#x?�t��P�����~���?L7�����Q�I(Բn�&zw�'\��4����O��;x��V�G; ~�?�8�O�X���� _{��B�SO=œOvm22Q��Ȯ�>F�$�ɵtZ�Q{�^` Zl��Q�M]�������N���0��er�f'FTD}��w~>����4�u0?�s�[ ��믳���_b��/�g���}�a�~��/~� Bd����K�&��v�(ϔ�=� 8j�6�#����H��b��b�^����P"�����JZ0b�TVM.�J���y~���p+J����g��;{�%R<�.��5�,��GqE����x�]�Г���c�1 S��w��߲����;���`3�ْ��)�.���	��B&���̚� &2���|:_=G�(��|/m�\F>���&����B0ОV�*�y|F�*�컌�?}���&��ښ��<s�L�P�\QO^�LLq)6��	��l��0�Ђ�r����x��y�B mF7,$�uY��#*Z��a�9��LP�"`�äǳ~���gM���y�~�I�&�_D��,���]`����{Pp.�{�M��rr,vx6��xθ&+ v�9�ոq��Ya��������B�+�'��Xu���h��)%�{1���t��jN�fQ2UG�L�'�"�7��OI��ӀA#�������@�s�@6�r?��@�讶>�M<v��s�����D���:N	���j�Yz`ZI�_C�ʋ��>lԁU�vݒ�!��354���y.@9��|�h����w)���D˗~�Y=M�Q���Z���U������k��b1(�8���j�hъ�m}��7�A�`Q���1�-0��Ȑ�K.I�'�Z�,��t(��Ď��������f`��O~����#�0��?b ���3�h x}�_Z!*���\W�S*Z�Î�B�Wp���N`� 9�v�L���n�İ8��x1DPǊh��B9��7�a����]w/��=��=�=�-���P�K�����1���$vK$�h��h"�t�㬷�t��`�R��]8���A���ߟg�tFb7esB�8�9��͝�믲3���z&;  �k�uA0E�[l��ؤ�z�����'m��w�2�]�a�.�������$��t�]u:(� �3�Mhcp	e��j�	Z�b1��[N>�E~o��Q���'��|;���TFY���Ę�4�?s��=�@h��U� S��16���x�@� 8A�������>~�\�VB��K/����cq.���(�@��Y���������_.��_q��)������}�g����TԮh�h@���{���
��BH�,B(����X�d�õ�;Eܐ+�`��n �� �yj�̺�)�@�����Z�\�?���v�x��<i,E�8�c�R�&�׿.gWϣ�:���	�n��~C1�_�{����>����_BpAD��E3�>�3ĉ��XY�Equ��
�~2g��'2��9|�%G�\�	�E��#����%�.=�K��m�����Ȁ6�����	��@�d���b$h��o(T�|��f���]!���\����y�C����O$�5�N %�֚iDO#H�4*�q�k;���KJ� $�;$�B�t�E�@��?!�4=?��#�W>��w��~;����?�1�eq�<�{�w HaW�����ڴi������T���x ��1�(&LH{��>�"�	�h<�	8���L9�98��-�]���s.B.�+D���u`�s�y���E�w4���!�0vM�:�,� ���
�t���	\u���'R4nq�^s����#�3(�?�r��������8�]z]��y���ϐaQ:uW�F4�p�iO�BU�d�}t#��ً6���� ����x��; '~YY~��;�` ��Zj�o�����27    IDAT�(���ƊFԾC7Z_���.+��0"|���߷O۝�u�t�xa ��I18
� @��M��c)�iUF�����uA�����y��ǩg�^�9#�hZ�׿���TPX��x�hh��^�S���c�� ȣ��,V��@����5cG��K ��\�7���6j�Е��5���of�4Y�s�-C�c�wh��E`����i��c��;�B"FmQ��ZN�;~��zVO��f���NЏLJ�$bI�s�.��#�Q )C��<^������b0�/]�2c//ڤ�� �sYGd|:G����~N�aQ��g??��mP�o����P=bm��
t�1�g癑�Y���89'�^U�ro�l����-j�b�0����!�9H��Q�<������˧X"ɉ��O={(͂�����Ř�P
�/솤��h�H�'5@р�����c� ��9@������y�^��c���`���7���� p�\�]Py�߇~�;�@
P�1c�a! �ʽ8��&�馛ҁ� g|�Pa�B�kKIP^Ai�3��#�7d�G���>��)Y$|C6�},hX\�N�+�K���E��}�$^�I�w�﹂��硔!���R��ԑ��d��~��?Ծ]g6�r��]��J��rTSU���s�EC�|�wI:8Ѿ�0"�� �3[�n�'��􀓟�l�d��X(L(�x�`� `�K�-�X�w�q�_�^�8�'&�cnJ�ʕ�i�ܷ�&���~���~;�Y=��mՒϛ��%܏z�(TG��Z/�Ȑ�H�J�ᢿ�cE;�/���>c��!T�ѷX�la=x�Hv�D�\ �C�@Rn�H������q<�����������<�'�P��*<_Q>����Ba1B;�o_\[E�p/����!��RAN�y�� Ա�by�[�v�W_}�89_vI�����F��kz'����sp��D-u��P���k)�qv[D�#�-�z"���ǞH�����s����<~P�w���ڎ�$��9��f��3;�Ocm�!�9�W��u�7I�늑�@��ud�\=ۮ�C��l�d[��~�cF��ɇM��p��l��2�!�xSL	��N��|ݗW�� b��DRɫ�k�Sgٲo��l5�=d%c�1*H�={��\]A�|�5UVE8�F���Ѐ��Ͽ�k����q � ��N:��W=�I4T�%:�b��X4` �5j11ax=�i���L�`��w5vH&���ջ7�
 ��~���.���i��;���ޡEc\Q����y�B������d`�Q]����?��ϋk'vH���(hY���C&���}�;p�0�"�0��XH$L��+�
	@�	H�*�7�<�&����)i�q��.�\V�*e/+�ѣ�҄	�ϓ�?�����~�~k�}ߗtB����� #�ҝaT@@ �E��8��1&�0Bt=���â��d�I��{-�W�V뭻��|���[��Mխ�y[��=�Ou������<���<�͟��T��FƊ6o�b�����X���I2�����=wr"�ց7Y���D,��zW���;�|���^�}_(��yԺ{{�g$Pd(��e�d�+�V�#&)zF<�����k^�j��h��3aae��3�Kֈ��8R鏍��:`���W���F(�`<=�i~29��F��UO�!T�x�N�d�h�\���(|3��Z�r��{�x��6R�K:���z�+(�E���qu���(a��r84�g���\t��y`>_�!��0G6Z�={\�%��G�eB���#�g������B���8�	��^�{�ġ��ݻ����QQ�0i���c��*<'J��SJ
�;4yNA�%��,�Q�<��r���;&B=�p�"dyw| r�J��u���p��5�o �չ��g�^�5�������`==��÷^�͛�{y�L��Ț�綶�V��P�YG�l���W�x��{9���fQ�4{
�~�w��<31/�(>Y��}2���ԟ�w��VB�5�f�:W*�-[�,�xa��T��*���l�����s{)�R���)�q3�f�@,�f������wO��'">���k�m"���m[��*L����X�`�KkU�c�a6/�	�S,�ȨdQ=���D�;^�[�z�N��ju��Y�~��^-Z�����y�sx����6:V�F�bfk׭��+����]ҙM��I�}��#"'\�C?���f2��į����#�F��ɣ�C���@D4��v]�M�0�c����;~��qo�q��C�&@
 ��ً�Z@])E�KX�S�XZ��}Շ�"�uP���(�1��@����n��5{�!͟5��A�4Ԑ�p3���<�G���z���|&a��y۹�^�-�(Y:Y��n��Z��iu�9���q��24Hi�X!����Ü������uA�l,s�k��f�w(a�;�B�e��((���n��;za�cHpO��:���6�4��������mOJ�6��ͥ�^��/���0]3%h�yX�t�z�+��>�D�N�:a<�]ג\���m���U��\�ȑv7á&��DGH��h��Ֆ����p|��Oʢ������n;3�P��\�;��2���}���6:ְF*��TճQ'R�Ǘ�T�̉F�ɘ�zPYߠq�b��`s6������Fи�����/|�A�Z��U>�s�\���ż��������)@���8v�r]���'��7�r�SWh��L����G�#�'a҇
QE�P*�wı�D;()KB�{f�S��¢�^��L�?Z+q�X�X���c�<����>���͋��7_w��_��V�^i54Vr*u�ow�g����~���y���˦)�@?�e��{������b��ɢ��p�ʅ!��S��#���ظ��x�����v�?|�P~��2Q���?�8͙�e�LچG��g����M��K��ƍW��;<�R��U��̳OM�8	:l��z�>�5���w*�_�4k��K읿�v��l�T�a}G{o�J�d�Lڵ���CL[�i�������y\ D� �4
�cҵQ �"I����w���hf����<9筷�;u�ی��H���;`8���q`�[�Ɩ/���|�����7��K^k��y]�	�Xiˊ�bnЖѬ���7�D�G;&��_ו������	�����?����^����-�ͺ����l��:d��r\�[
�h�0��A(.c�x@|�3���'����J
��p��1�x������c	��@���IL�
�M���� ?�O�u�[V��T3���<q�>���5sI%�Z��nW��F/�ݺuvͳ��|�l���dl%��C�8ξ��x~���?��I����eng��f�XC�x�T@ɲc~8�d�ŋ8M{��I{��'m�L��ǜV�g۬X�x�E�����l��%�\����V�Xa�Q�X���i�={�xhh�����dO|��׿��v�O]���~;u�=�k�ϟ�S'�˲�H�ldp���Z笥����c�S�cO��dN���N1�_~4�OZ���:�)�3���#g-�L[&�a==��U��86��&������ݏ-�Ϙ@��1�R��B�㌖̢��������LlEca��b9��7{��; �X�YE-���͋�G��x�?�2�gh�>�`��gº����7���;o������ODٽ�i�7k�����)18�y^����ONe'#9�6 �� �!G�
����B�`)�
�F� ��/��K��M��ۮ�-�iX�D+G�ի7ؚ��Xjxm�l6�a�����yFm���(l�&Nw��F�}"m��G졇�^����J@맪't��uyn�
�U�kTG��w�����J�UR�V-��[�a6^(��c�v����7���$��_��_��u�Ȣf�'.�v�����/6��O|���=�������&����Ä��}���|�b�U��o��/m붫lt����?�ٰ,5AJ劝<~ʆF+6p�lo��o�9@�Z99O�c�������R�?��Y�<f�d�Μ9b�=k��l��Y��?mc�����������㣈*7���`��%rg��s P6'��E3f�J�D��QCu�K��ht<�?�g���#��2��ٖ�[=�h�O�s��#��ޫp�2��١c�����J�'|O��BOhМ�c�	*JH�� @IF���}�"@H�C  ����]@(@��	T��8��|��O*Y��������K�Imݚ�m���,���*�`=_B8�;:]��5�8|Q* ��z�(��o}���X;U�|G()��k��<��J���=k�ʈ5�e�;�g��H,sK2�fǏ��b�aǎ�[��N۾�j��=��<H�G��d�ό�[���������J��{����ۿ�V�n�j�?�h�]���"���b1r �r����<6`��,;|d�6l��)Z%� ڀI��Y3�ACCӜULG��^�÷2^���\�a=={���V#q(�m��� �i�B�2�>�l��e�F�9��h�܌;>8ru�b���,B�(@���d�Q=�lp�)�+ |��;��/��"��=�:B�G����@�a]P3�?4�# �5Ƚ h-B1�.��8�cD9�
e��\�*�rh�q�����p�N���`9p}�'h�XXD�`A�(�(i��fM��B����i��E�D����\�m�Ԯ޵���%��m�u�Zd�_q�Y��J���HeL��'�X�Fl|�>���@1����o���Zd��Ԕ"� _!����c8~h�����l�ڥN=��+ǭ���}
�Z���=쾉ѱ��Z�����wXG�l;yj��z��S��[v�ghx�C�4Қ�+�W?�^/��ݳ���7��y�c�{�4N(5M�mhpغ�{�����c[�&�I�X���h�T=#��DLl68q�ԅ<�ٜ���p���IT=sq�8lgN���[+�[ �筯�k�����sV_ �_�3o��4'8{���Q�)�q%�B�=�*����P. ��������誉
�g� ��C�q�j�ε8O�;�& .JJ�E�9�/�%�&��r�u��T�kI �x�St���C�����uT��5۸����|3��KY�e\�#
�$,a�PO�8��������_*[.�r�/��յҮܴ�2�v��	�C@5��8~|rQ����sv�0A�1��94|�֔2���r�X "ð��������|�6o�`����w����b���B�n�=w�2��v��/7�S�|�
��7R����۩��x����u�݃�C�>��=�6�j����T�f���}��u����^�����6>Vp��d�l���9r�R�Y����bӎ	�gS�� W����H�4�8�S�Ntc�l�yq����D�j'���=�X�FB���Ȓ = ���z���J���X�("�y15-�8z��[�x�d2���_߻�4Τ�,��TV�����k�������Щ�s���y�����M��Rք�		��1���ֈ�wx|�<�YϦ���u�q�[���Tb�����*߅��`_�g:���/Xow�����l��Wx��<�u������k�o���h�r۵�Z��Ky�Wwx{;Ԇ�������D� ������U�ư�H�D��̄�B��88�}��_�(�9sf��C�}L�wTm߾nK����Q+V������jG�#�K�qԺ����En���}�|bhh�7��=&���������w��_����~�N8}�J�b�O��P,ّ��66^���5��ҫܳ���I6�q��MQl/�+���(,���*��'~�^�h��>���O=lgΞ�������:M�H[6�n}GO۷�����,��l���d�ǛX\<�o3� (�T���&i��p	����څ]\"A�^��N�y�ֵqB�-v�K�I�&���h�uX��.V�tr��}	E�85F�v���,l���8��^=ח�YA�r��zg:p��y���m�%�b���'�k���C͈���ވ���uA���n	+Z�Z�(�T��͌U�)�5�~��W[��o�6+�	���x\����#�4�^4���}L�oYc8�J×D>�|'�D�#�����)����b��-����?y̪��[��2/�O&�e�N���K���?d��s���1�����+�_�p��fjI����gQΞ�i�|��l��%�ޖ���_�+�Z�6�_L?�;��Œ�����Ƭ�t����w�㌍I�6&E����LD �S�� ���jT�W+��h�,sm�<qB�9`'Ou��\)xUO�Rx/��}z�>i��,7:�f�r��?tBJR���M���P|����Pb!�zC�V@h;��&�^Cm\�ǉ+�Ix~��f�s��4��u�P#��s����9�/IJ���P�,�����	�PP��-�f�L�j(�4�\;l��K��b��Y�{����3~��8�{����|.e�zɮ�b��ܹ�s`���wȵ�{M���k	[�z�U=�&�}/��I|��>g��/����;��N{�k~ƅyDt1O�����N��O��r�>��}�ha��S	;5pʊ�1�1� �z����q������7~�k](}��G=˻T�|�/��$���w����Ї'���j%�F�[n�����6V�F�h���sV��G!X4s��e��6tn�N��5Kvٛ�����<B�T��E ȓ~Ы�
�:�Y({���I$B�	gQ���*�P��>Lzil�Ν;c�:����Y:8�̒�W��И������k����k�y�8�E�}BS?����� �ٔ5GY��k~*�����E�7�����e�:�����t�/KA>	���-�
QNa$����)ԶC�Z,�@W���JX{du�,�4���JP7[*/U�!�/��kVZ�&�?��7��O9�R�9]Y�;���uG�xT�����Ȗ�x�t�KĹ�X |::���@�D��������O��!��R����������ر�����;2|�
�v�d���7Jʹ��:�y�IK����s{�E�?�V[�d������w����po�
b�^�ɝ�n�����M	���Ă^�|���]�b�ͷbaԆG��#�|����D#2)�eʽ���c��̳k����L2�rl Ջ�!�VzQ�S<p�lZ8B��r�h���6�&����5��g��=K'1�Փ��|QS�0�k��B�H�Y�v�z3��	���"!.�� ���7���4�f�#&ː��<iѡ�>ḇ�G ;-���}�Ly����.��9�C/C�<�eB���Ofq�<�q�Ӹ���BJ(����T�<%��f�n�g�Q�����-�({�Wi|��u5�Q�e"��b�b�sl��^�'s���p$����V-����)��p�b1�Z���C6:%�(#��(!�����[�*6p��>t�N�������6K4�^_��Jf슍[l��U^���@�,�p�M6v�Fc��h�x��TEB\�u�ַ���Fm��.;sf���N�BR�}�Nۺ}�D��K�B���u�?� p|�m���P/��<0�	�ęL($Rǽ�b*��'�}�8���Þ^�j�ly��b��6^�������M ��������{��Es�����oH?4[�=�/� i�D�6-�?3QP:Oc��!@���|�eYH��y�V��]�#��� Y�u��K��*,�&�3�4����v+������m����L����E�H@�X����,YBmh��F��XH�@�.��a����z�T��W�	��I�ܰ�J��[�yKPJ�����w�    IDATa�1�>0p�>��>g�Ҹ+R�Qf�*�K�w%��P���	�ݳ�+�
֖�X__�=���=4���âF�+V���o���̙��B�9��E9tz��gF��n������_�J�WU�Z��Y,�{ӊ��Fn���I;E�0o�Y���p����=���Q�(&���:���P%,TZ�7����T��@�ؖ���5m6ɲ 8@ǿ�~�N��X��=q{:�p���{���=f�c��f�^%��[�bu$$�+�x�>���GH��+c�����;�R���m�N%<D{|��K���t/Γ�PXg���<��s��9�<r�N��J
�yo�y�B���C��g���ZD )�?�~B�*O�
?�'�����][�P��7P��J�D��U��j�T#�?����Ջ�}�e��͖�G�I���w(������1��"�oo���>h�����y�����w� ����16�C�w�hb?��
7V�U��`���J�IgG�G���%'%0%�����xN�9h�o~���v,��%�Qѹ�>3�o�s���{%�D����.�ȭ[7{���~����{z�%HĿ>���.��nB�S-5�&,�E� `A�!J�Ϳ{��y�E�ڏ��T~tޟ�rq@�U���,۾��@�/�z�liZ?&���s��i���R�膜7���K�)�-.nIg9 
9cƀM�u���D?1��Y�*Q�xJ �2��/ R�fb��p"��P�G`c�q<�AT�^c����9��p׆� #ƞg&v���]�~d��X(�D�l5�x�,lz	M6� �g�W�%����[��{�X��D�����pMţ��Y��	���?W���M%
��g,�G�J��%ͼqnX�q$�AIz/]������	O�"ڇz��,А�y^}�&+Ǽ��$v5��'i�5{�]�e�G Q�n^hހ?-�3������w���ٟ?��M���\@��G���}����Ԍ��E����[}	%oԫ�k˻J��7�I%��D}��oG�qw�tTl���,����i��1������+lێ�v�����Ʉ�g�r`ч�t���A�%ٚ$uQ3���L���OD��6��#����[5s����#�m�T��k%��F-���B Q���}}�v���c�굤�]�>���{�.�CI[�j1�� �f �qz!`�v�V$)������a���G13	U�Yuo(�FF%�qŜ�: !ay��l<
�~+͘��l	��������͍�M���4�H ��zTڤ\��}�A�l\(��F.�$�OB��|��'�G�Y�Ō�Z6�.܃�PuX�EX�=nٲş�h
"@�*V$�+�'������Qh��'�źe�B?��Bk�8� Y`<Ϗ��5�j��U�P�0�{'�����&�.��	���Q=���m��N����^�皫7��)ژNd�TnX�m���3w�OC��:��6��j�Q����g����w�����n��V��#ܓcM�?B����߉R�>q�w���Q�Q@j'��")���ɧ��y@�Jd��]��'��L�󟺼CӨi@e�+CVC�c1���dܵxMJ=������I�' P��?�A��{|)S� �0Z�����j���9}�z?g�҈�57sm]v��xTۇ�΀������3/ry�K���j	���Q@���#��	�c��ËEŘQs���%@�	� 4(�����E�y��G�MŘ�`G���G  Ҙ�gxX
�Q����� U�m�|��ا?�ihr4e">���fF � P9���F+$������^]��C  Y�J�`� ̈�WD�.��@E��]��A�I,�Y#�1`iV����r8l��y#f��C�I�����Ġ&e#�;�G�ERm���<�04ɅX-���� ��$�"��*��9����g��zz[6ٰjm̶m��v��̊��FK-a�L���Zn�6l��IZ��Jw�jO�?<;�V�
��}�3 P1o{���C�kpg<QX(�G�&(�ЂcND)�*7�NtR@O�'�1�¨�h��o�u�g���?�#Gd���Z��u՛9_E�4K_-��-@`�g�e��� h��[����W�j�d]�.��������iTk^ҹ��ɉ�nQ3�FT������.3� '�ECcs��Y��� �G?�Q{�k^��-��L�� F�B[D@0/l@�z��Z�	Z�� 	@��Jm ��4rd����c4��kM�b�U���<� �l� �(�v-.B:g>@(����;k�͏@C�N�0@���Z@�G���'
�!T~4��ތ-��&H��d]!����ð`X�|�*���I_c��cҌ	sûBePH��5<7�KDy��"4��v�!�0@h�>܏�X�|Tj�#'���J:������@TϿ��r)�re�vn�ܶo��C����<.���XǬ�6>^�j\ٓ`	�ѕ�j9�ԫ^6����
���}�{<��g�b	a��֩�
�KM	X�5s�5��q�~���w�5�x�}Z,�j���XͿeU�x�B���P (��9�Z1�!'�̿q�����j���aΫQ�%�ܻ�����e��O����Nؓ������rVk�����#66vk��bY�����{�}������VҏLd�l��y�&
�r���D��� � ���1��$�Q�8x�cs"\��;�U?y>,1�h�9�ȓ���Ei�*;V����$n\��h� *-3P�� k �x���������]w�����@�g=�BQ	"@��L�6M�i����]ԑ�5� f���tPj\���E�	���L l�������a�b��bC��@�1N���xƇ���ȉ�����'̎n�W�6О]�$�����L\�?�ߊ����k��+��}�Wk�^j+�\i�:%*���4�N����LD�`&�t�A<V(x�^��GuPذ:��+S�RZ{�#��X(B4��/֏�����G2�5�[v�~Q�\����hIi�k���P�H�7��\
�G��;�1�, ���%��l��ג�M�^AC�ٹ���'�F�>�ԸOؑ�1��MN3��zRҙ���3�p����d��w��0XGP2l*U�d�Uvm ��PѪ��DB�;>|  ;�8�0�k3)���C@��riV�g��M-M�gCp��w�s�� �?��s"��]3��n���~Ο��������D���Y�\��P\��<��E�@��z��"� ��yg���̀���JQG_,,31��5�c�b�7��1�Z���`e�<ļ3�h�X#<��1Y9��J�\ɩ�B���������|�T;�k�F۾�rK����9��z�[��*�6�V�'�A��Z�����#~�<�b���r�|�9ғ���wG�S_|ƞ�fܨ.���|�~��0�K�-�I��!� ��hi����o1N����wF�����#��T!�#�r���Q6���ߘI�\hQ*��h��X
��h���k��7,�6;kǎ����yR�s����3�?�����������F� � ��)9 d��!�D�������C�x @�#xo��c��E�b̠'�ș b +� ;ԉ����� XC�\_�	�q�H�h68���������@��9~�"���t܃ka)��o�[����g�Fk�Fh��:2�� �j��
Nj��x���NW�AG��}�N�O�ϸpm			F���X.�(��@���c2�|x&(N,+Q��������&�d*Z�����q��1���*�^<����F�*6�R[�f�͞���;$29KT�zD�e,��ɦ]������>_�zT���c��T�9U�g�{	נhq�a��K�F0�\Kʢ"�Z�����n���}n�whh�=Sq�tih��Zf��t�Ĥ9M5��|Y ���hB�)'����A��7��ꓨZ�6j��!;s昝8�cV�!�_	�Kz��Ѩ���>4��G������@�KfY; �$�V\04`�JX�M7��9�GÇfPC�8�~E��^6��0�8�c�9�s�����8D���<#߳�)ԇ6�?�v��X�Zͩ�	x�ݰj��p�h�8����K�X��@ A�`=�}�4d=���7�e�@s�R �yg�1��yXT�3�$~���&4 ŸBc��2�9��	�*����!|��4R�C� �emx�z��~48q����2�p✃pVn��k̉O�S���9��Ba7���{���Q+�V����d�ƸY��c�,a��$;q��<���ͷy�;��h�T����;�z�h���P*<4�ֻ��Q�G�:o�@	;�£C�AX���J9l43W�e����{*�,���w�Tܿ��Pp��C�˹����5YD���s4$L~�^���0KT���G�T�eSu��j�&���NB=�����oT�?k��<� ������4PQ5
d18E����� Z'�1c�E�3�aB�) 8R����	x"Դ]4���
d���V���������w<�V�/4�k��b�p=��`m�vۻ��?BI B�{Q����Hy�6c�?�*�8[�l�J��G0����;����F���?A�T���gM3X<�/��cqM���r,ϧh"�Hh�r�ù�0h$�3��
���'��O3��[OOTҹn�y�Z����I��`Z&=�GJ6g�����a)��I���l��g\	#��λ��9ͷS!7:��yY�
"�~������؇�������l���-Xxیl�8�K�ntw�0�q�prB�j�2Y^2��[��8�l<b���h�o�bO?y�x�?qι4�a�nƶ��0���o����ڻl�P����g)�����S	.Z�DHP�Q22��R�o���3����^�"���dI�����cj-M��C�h��+sqmy9�B�D@������~���uq�P*PC�,��D!�y��XD� ����=Ѥ�%ᫌ�Ve�� �;��b�f�xVU��$r=��wFH��ܛkb0g֢��/���a�w#��5˹ⶹ&τ��傠��X��"��S!C���/њ��D�Oe��/Xo�a��?:v֮�z���S�l�0�;�L֪��n�:V�,���WY*M[Ժ��qͭ{�{��G�c��Oi��eh���B!�5�R�C�����R_g�
��֘07��ߕ��
[�y+����U`�s��ܥ}6[�'��,*�k��Z��1���N����A� �w����W-Q/��fuം�,�b%K1��ځ���Ǟ����'}���r����b5s�F�C�$�Yc	8C�����@���Q�ތ!�E�	�7��ax�"M�0И���$ņ|� ж�x�T�.�A̛�6�^f;@Z#<a|j̃���%�Z� �ϵe١y�
�û���������]є��.PK\ޝwCx�[ ��&?m+�֋�5�D�qo�K�1�r@h��:NYuSh��W�.�$j�ga�3P]�{��	�����Ԯ����=�MĚ�y�5� Z�w�*��^�vݼ�&8��+⪞�"9|)��qGj���M�m��+,��z�o�ޒtK���Za�dU/�\�|[�;~=�2���pl�+|��&ٓ<���\�Q�F�	�sQcr��]�5\g���p�$E�_�F�Z���,\����җ��������i��3�,X����Z�)TO&1�b�i*�xX��X��o�y�%幷��l��Bi6�j���h��IFo٪%
WQ�6�`_�elp�`�D�ʕ�,q�˗-�����0�a.tލ�6?!��s -�b��@	`@q��Frt�'����� T�7 e�����+�G<`�#�EH	\4�2�����hL9^��O���1�z�C[���%�U���yމw D�l~�#�����>Pp�D��`�6M�)`������P.��揟 ��Z�̬]�%|%aƅq@�p<�
M�{a����0��<B�s�P�^�R���A�u�_~Q'-@��\<�g�
/�|��D��Mٓ��kE��H��Ymf����)����@�'V�&��HY���\�͊�(@�8>�}F%�P�%ӕ����(2֒
���Pȅ�(�kM��0��f�*��Y����o��o�����ӄzJ"��*�]��f`s�  �]Z�jvȡ�w �4���S�!�P�tp�:F�)a�`���CV),�m�yu�(EͿTI�h�j����3:-_F���.nw9
%д	xW���`C! T�5 ��ln~'�@�)��#��i�r�|4t�08�*<6�~� x.�A~��&����>D�i��W+B-\�7�E�p}�(izh��MJ�뉱A;�U�F�O<�:�j�+34
�B!��/��%�9Z������� 0��DQpO��\0'�cM2����X�#Qb��S~"�p8�ySY
���r�<>#�V Z��h.�d� �~X4��XOO�u�wX�4b�d��U�4<J[��h���g�Ξ��6n�f	�zE���1��eU/��"n�駟}��|ܰڇg�0�����1d����h3�Z�̍���a����1dO�\�l�߳珇�o���+�����ĝ�Q�d^n�^���t%"�́F��l��
ȧ�Ρ���-\2��*ɋ�'��������Z��Z�D լAU�l����g��R#�n�/Yk+�/���HR��q�Ffч�Ei��5#�_��4om
EN��F����Fi�:�ߡ(�#E\pOi[�V�����

-/��d��y|�dѦ���ϵ���s�4QMat����QD��$�Bk��d���T�A��,S���hL�!ϫ,w���3+��Q��9��q_�%��k��Ƶ5��;O�o.�����cL�8�S���s˹�(چu���K�X�:�e��(y��i��;��x�n�V�}��N_�"h�h|3n�}�'#|h4\@Wc+k�C��;�
�C9\�1W=)�%�f�0D`C���A("4�(7~�20�OD{
���Ok���f0����%����:�� *�y4=8LņK L�
56�xa��{�c!���I&jv��S6����esIKԫ��ʣ-:���}灇md���x������5��bT�x்.��ؠŰ��=���yKi�l,�IZNH�79w%�Gi�y���X���ϩ�' �Uǵ��#%ABBڜ�Eq�l��tM"kI� DJ�~���7O���Z���9�g���y<oi��IWֹ�+t�A�r@r��Y'��X1ךC�'Q������ʟZ�Mt��:]�l&a�ڸ��v��tnT"���m�7��-�=�����:w�9��Yq�lt�i�Ko��;~�-���7�4AI���� 1���"k�c�
&V"V��=QG�&(�'(B�>�Kx%`*v�e�o��3	�+76��8��Xf��&4�"M�c�˄�z��8��H��{Q"'ؼd�NI�$��w�#6<|��U4\VQ�p����a����~�
cKg��J8��{��b���N�"�i�r�3C8��j৸T��j�(|�kl�fB�I�� �����p=6����k���mq���G�&��E �@��8_Z��$��>�X��:N�������B@E��}��r_{�IK0!Ƞĸ�4x����(���}=C(�$����$���CKq* �{Pҹ^����aˤ���!�r�z۹�*K6"��)�\�P��l��e�e�.+V�6,��{�&���F�-�?���>h���֬��N�=e������C �J�#c�>Ƿ���^�Z��QLQ4�����/�����>��>�B�>7���v㍯�&<I)�aw>���޼����_h[�l��wy��5�IDy`�� e*����A��c( �*ԓ�t�3v��a;}����/    IDATU�c���(���\~����?e�Σ�Б)�&��K�{}.V��(i���%8F��%zi�i��t!�0�3��K�4���e���I[�!(�u�*�%���s�kB�c�f,����OBCt����9*�gܸ�'�{*��"ǤK��K )�M�U�c��)�� ��Ѹs=	EJ5BY`�B~ 	E�I��&�?/ ������D�oV�M�а7Z&E�fT\.��]�,�d�lպKl���f��&b��'
�������OM�d(�K��d,�ې�Cd��Y��ɾｷ[[[��mY/�|��q{�{߷����o`Ū��;���a�t���Pw�����o�/h�/�����S��K�w���p�l�D�������Ν0h��� �U��⥫�k^i��Q�)�q�L��~E���ӂ���Q{<9�ظ�>��V��&�����f�L�Ϟ�Ç��b��k�C�g+9v���S���;ԓI^5����o^��¢;H��Zn��n|��@Z&?�'p�w�G�d�:�j����- ����F`���l��d�9N���Ӑ��=��7�D\O�o��hQ$�^xvmx	{i�>F��k~�ֈ�AE�	h$T[�~j���� ��.�z&���%�{zڧT�m[/��;6y���r�b�d�.{�.�5w�e3m��ztl�#���z�j5��l�C���Oz�s�LFY�a���5�ߎ+B]�Xw�2BUٕ+�Y�R�Ju�~���l���V��-�H�u��>�.�|�m�~��)A�L�����O#k�g �V��=����F�x	�¼��֭o��
�C66|�N���޽6Vt�ϻ��='�v����+I�;o����q��r�<�f$�[���Ą��O#
ca�
 Ĉ��*�� �Q:e����ؑ笧�+���\&c�|�uw������6�sA& ��F�L�A�����H��}fuF��DE���V�(c#�(cE�	ILQ��W�6E8'@U�i��[�7	ݛ���*��n���s ��Һe��9
r�[�{Y���k&�ώӏ1����y�$넱iV�uC��z���Um�����q�'r���m���M��b�F�/]mk.�ʒ�v+V�^�'�J{/���X�)K�纎2��Iu|�Ɍ;g�KE��z�����{���g���;�����ș�G��{�<�φG�hR��
R���F+���]��M��	+���hѾ�կ{QH��~�VY�/gny��J:k�9O�_�h���i��?��-Y:���<u��e4����ㅪ=�o��������.�p���夝J��-��c��6�8T�>$<v-7w#m�T�����Hة�����,����$g�ݪ��&x~a7�FKs�����'~��S*VX��ЎD��8�\T�����U�� watl������Bg��q�lB2Y	uĤ�C$���$�!JK�ҶC��{`��k���;D�8%�qo���x��Y�8p��O�h�ٯL�� �N�	��O���d.�?Ɓ�2j"ϼ�S�p�a��/O�U�|�R�Nh�����?��zy��;7Z>mV$,�Ҷ᲍�pɥ��tZ�R��D�9���9���s�t2�@Nm'������=���y�X(z	�H��LrY���?�����z�F�O��O���Ҹ;���Kh����6pf�j������b��^����}��H�iB�_�I�t�\�of�aK/�z%��R���'v�+��$M�{�[�i����cG��V����C�e�.O>Bsd�PGF&�f�_��8[4?�<�Wm�B��>��U+	�fR�˖���C���I�T�L۱���f./,��O���0�����O ��fc�H�v-���������C����p�#:I �Xq��0����>e�)����x^�&d]s�� �ʼV�l�"2b���z>6*N8������%�9aA"�W6̝�"	LDl��u��I��Z��#��x���A[�j�+!X'T�Ĺ��#������Ci�G4�L�LK����C3�-�.�]�l�|�zѬZ��K����vX:�?8��Rz��>$|�͒Q ��4��mDh�];=�\�H�#Ɏ5E2�Ah������.��w����_�����C����s>�POc����{�::�ّ��v�ƭ�����^��pw����:u©ח5�Iv�-{��l�X�W<Bf�ʕ�[��[�j��ࡽ��w��j�g�8��&�D=i�#E;q���>=G���;<}���Ԣ�
�(��d����pO��� A{�yal-�z��&��l�'{��@��=s܋Y	Eu�W�OU����1���S�S��r˥���Xp���h9�È�j6象<���pp��.�(�' ��LZ���'��0��"��|
��tE�.��JHK�秢v�`��D5���`�����/x6�9��<6w��-A��P�L��\_���A����~e"�MO$��:�*�#~r�>ƃ���ь�������j�yrc\Փ6�1��s	��kǕv�5��j��UzZ����m��E���T�?�ō[-f#'>%! tJ�D4e5Ŝ��F�&un#󙪬R�Kb�c��.�?5��Wl��ˬ���{�.���3Y2���S,�j��g�-����;u��M�pj���!�
�̥}��d�F�%[�z�}���3�(��O����W_����w�5��d"c�C;v�U*i�>�?Z��o��J��|���J3FC����/�뿣ɲ��rQw��k�^.���3���g���&�!��N�[w�@Tҹ���Z�Z�}�����Lg"39t���+����dI�h�	GlowNt��elr�)�S� L�LS�js��M��B�@��	L������|<;N;@\8s��]Ř�;����u�������Z|8��9�g���|hͷB?�t��Vu=5�x'��8`��6

�$�D� "N���-���pή��*۱s���-���IZ��0Kϲ��V���Kl����9&��F"�0S	s�k4�.ؙk����	س~Y��]��Z�R@�,��s���y���X.��cǎ����HФ�ܡ�G����ђ}��`���V��Mh���
��8c�8NG��,��d�:�������u��/~���~��2;ܽ��Q�=��C�#v��	�V3�w|Զn��5 �^�E#'��@���h������{7'�ςB�g���� ��M�$��lh�%%�g^��z$��������X�Ƒ�nk��ˋ����
� J}�G�$�86�\��X8/��:G�XDu�0�Rܚ���<�� :�%���c<�7?
J�P��&��͇&L������A�����q��=T���/D8V��!U'+�9���ޔ��܇�D$�p9�~Rl�|#����(�-�$�Ph���z��Λ�q�;
��}�9��7�у��
�]�H��
��$jhZڇ�==n��#v��+lێ+�Ny�l5/�l�U�d���]`۶�Z�J�9�T�lg�J���|��]wOXz�e�4��p��)�֨ΊR��l�)|Sp�(}}{��o�/��ʵ.zz��Z�!�����Xɞ}%`����Y���5��5�N��v������T�`����f.�3|�!��-g����ys�X�������֯_i�cC6<�OF�����;f����l�n~ÿuPB�S
�pO@�C��P,V��͌_Gi�L.jD.���E��M�qPKT���'�H�~k�S�d�3}]�E�I�[O7���9�����Y��<_��W-�kw�zʣi�_�-Y��n�G&Q|7��MC���p���h'~2n}��@��]�M!�F�6 ,�	�Bgr�+�J4WsC.�6s#*Fs�d(9�$�(d��z:j���J��C�b�K����8yk���߻��.�8ʹ�����.�}>@��%��`�'�7�}��1��_�mۖKm�+<�'A�;B=3yk��l�P�9�ث^�+)~����~b�� ��wMT��C2( ��)�>�$��K��`�}�"a�(
��=��7��3ms�̲��38m��y���#�ldt��O���ڛ�g^{�7�yv�>/��E,+�e�o�
�U�L��J���M7��n���f��k�#�$h�,K�?[�9WΟ�S�m���������S>�Z`�q�UE8A�
y9���'��aѱ8�j[��U+E�7��P�8bV/Fez)��ى���s�mx��>�锭\�ܖ-_9�����_�� ��r�~�~�ߏŷ|�R���W��Lԯ��"�І� �z~�w~�#��}����&���f�`m�	�6�h� +?Q>h�,|��\���&��1/8e��XlR����1�jnx6Υ.��k hb|$4$,ࢱ��D��I��d��q�a����PH�Ї�}�O�����w�r5xq+%Vx?�k��1�k�߈�Q<7�w�>����V�h�t�๰4�o���PP�;���M�>�a�C�#Ը?����Z
��x�� ʵ'�L�v���lTҙz�����_��.�b�7=�륚�sY+��R���ZmX�FV��Q �RX8��t
�>N�5���N�@7���ظ+����cL3醝���s'm��Y�JH������1��=f#�{ǯ���`����}��}Oa�Lc�-X��/���|�L��9u'�F�J�Zd��Kv���/���6����s��SO��J�FTK"E�� �,�]���;V�dTT���Z�1�p���lf���" �=�7��b8�y�RqI�L1���U\@5j�*{�?B�\%3��,w����96^"d�b��|��X��
�޴���}b�R�ģ~�	���t�Zf��t����h��i�X�� �u����ȣ�� (m@J��!c��� 8����В�3�X���&��y�&>;Pо8_t�TH�iL��9<#�}�K_�,����0f�a9`��� �`��B@vZ.�l��=�Ԧ�	�L	`ʈ`Ma8��J�v��: J�φ�2�D�!�yg������.X���˚�3�Y�Șk��z�|x�3���5��FR��Nh#��yg�@�E��q
�yE��T�a�^��d����d�$�����V�|J2ac�g-�M[��4��z"��(K��-�J�*�/{�$<q��dv��T����xG�Sy:�8S�R�(41�˹0d�iPT��[W{�|�z���(�uKeӖMe�\%���i۸y��[{�c4�_�K�7���Tz��;s�����}ph�]2��xs��HZ%n�<>:�����z{���R������������������a�V��׾�&K��zł����U'���bƹ�4���'N�t�s�� :6��<�q�8M��mu�?q܎�v�?�%��:��L��600l�t���B�
��X��J��:c+�'��;�t$!pQ�����fuL4� \٬$_1ԭ��"d�D��%2�1@�ط�9S(>*��;0�h4"���k<_���ƕ1Ҹ�a��3��x�d��0[��b�)�E�C��*j&`I�c�I`�d/4Hx`@��[h�p�1T�7���������h��8����XB����.�hu�s�?����ܯ",5y8�G��p-|Mh�{� `�����u m�lƁ�&8l� jd4Z�\�5�����>��D�0F��%P憹b-  ����IP������V}��k�9s;�R������V'E��t�=�6o�f�k�v�Xs)��	�60?�G>�)�(�x�b����%HY袁yO�x�޵Ò����{�g�'�ǎۙsg<�c��Ev٥���l��n��Dʾ�������}��E=^�IF`:����|AΛ=+���|s]w�5�������>�4�����uk-QoX�3~�644�?4�o��f��h�y�r�ı���h"^����ب��	��ھ瞴3T�L�,��Y�R�Q���t��C'�������^��s�-[���5#��Bm������,b�n"�`D''�l��e3�b����Ip��Izcs#h ����3O=�&36r��9��	P#�µxv	�x������2��46-V
�E�/Z4��D�V�GQ�G�]�[�/�����y��Ra�� �x���&ƀ����# T�z�k@��X^��>�4��LX_<'�������1h����'?� @#��C�@� �8�Ʉv��������Zg�c�Ag�8?� gm�[�_��`�P��(@�o|��'�SZE�fj����P��>�4���2|�N�@��֟���x��/Xb7��j#i��:���eg|[<t&���½h�B�19�qd3��#ㄦ��\'�(w�wݾu��!��(<pp�����  W�Zg�]�622f�]�큇h��W~�H�L�3��۪�{�0�h"Ж	�$������WU�^6��ѱ1���v���kAl��,Jܒ��F�q|��؀���������`)@�xDJKͿb��>j���d��5~*�B��l��=���=aC�t����YV����ޭ48����Dҙ��>���'lvx�
`ġ���O�k_�:s���׿�5��W^���F������.n���ccqc(�l,
�b�� ���>�FT�]���VZ/�B�)�/�e�h]���Q��SҘ�8t?~z</c�,nE��,<?�����C <�ll| Dƒ{2�h��?����k ё�aJ��̀P�3�!<?���&c�u��6�;� J����F9��`y�����8Xdj􂠅��:P�Xm����{� ?]�L������"�Zh���t_j_U��^����Y&I^J�Ն%3Y�d�FƊ6{�|���<0�.x(:XfШ�?�K��p_�v�ڭ�[@�yG��S�>���������׽��8j���A��j7�(a�"s�\�H��������w��Q$*�MHw�O��(�\🦍#`Ƅ���h���h�L�Wl�-���Ƥ�_D�@E� �*�M���j`�"�p�hЄ=)a���Xm~�v��ΗҎqJڧbGz���'���4�Q�!w�&��p�){��O��%�;�Z��V�p�GV�T�?�@ |�cI{g��n�J���=������G�,Z;|�-������Zԓ�?1�)��q��c P�u@T%m�t�����"���wm8�ņ��A�0�r��@��.aYO�<��q�D�@�BQ>ʁ�'�O�K�s \z�AK���|���s�m���#��oG��G�=���Z�ǃ����f�l�a��5�X�PwX�� �h���g�0( �\���u�څ�йV�� �=��P�Ϛ�jb,v��I�'��xX>Z��͍����f��;��{�r٤U��z�z۱k�%�eW�Ru =m�ɜG�\�y�ժIKeڼZ�C����G���}��_�E��G>2��b|�g,w���*ժ��,T栽c�]q�+�b^�v��x��G�`V�Ç{���r
S��N�
��gl��t�>��,2@�	Ne��F�*e�1Z8v���j�}#��бǩK��Y���9j "�z�$XR��?Q�BB%�[q����lxp�FGO���i�}(E��s�Ġ}�[߷ᡒ�ۢ"j ��UK]�F�i��cݐ�Ef#-���/~8e�Xo_�or4B4M VM�т�� 6���骫� �	�-	m<�m��;(��h�|�8��8��^e���f���]������N�7�6�W%P��`g�a�+GA�E�T\�(#9|�;�׀��g�~�%�)*��b�������}��|:
c	��Ppli<*�O
��u�������r����sq_���ZQ�@�J���zrT+(��eMqM��g�r��8^TG���O��Zͽ~j>� ��)3|[��v�����
۱sS��e\#�?a]]�mΜ%��5�/Yn�z����?�L�ӗ+��>�G���E@~�w����)J C�bY����)6R��1    IDAT�gfnU�;��f�%B�#b�����K/qg��X��A7��SKD��{ǭWy&/:���?s���;��/Ȓ����'���ظ�e�У�^�s/��p
K)Ւ4���b6�������ܤ~�m��T��tf!Q�`J�oDF_[&�)�=m�O1_'���#>n?�d��H[�T�K.Ygk�E叧4�X�{ m���F�n�3.�0��~�X�[Ex�A�Y�߷ϳzh9,l�� F@���G����E�1D}��|������A�I!P,a�Q	�ph> j�N,5Ȁ�����>����.�ڝ|xfq���tM����a�����W�ʩ-��+?s� exVh�2��zr����"����uO�����&|P�z��»�""�k=N����h}��� <�ƃ}��%�����; ��<�s4��/^Ѥ���h���)+m˖vݵ���;!��x�ƆKw��+�^��;��A���{�tųR܍����r�{��`3� (���r�χ��KOF9@h��e�q~'�8B���3I�����"��C��7�֚d�f.��t�Ʋ4�x�ġ�?��g�b�4C���D9hCiSPd�@5@6/+��s�펅%z�Ο�:U��H#JZ:��.^�D���{��g��+Ke�Xo�I{��ld���Od@�l�b��}����X;:�"!��c����B��[�0�<!nJ�
5}Ox�{Ȇ�����������T�V�-����t�{7PÇ�P����59_�V������\�MO�)`h*��s��
 6�j&XQE����_�U6�m��6��::8Xq,����/��}�����d��<q�>��(×���d�9j�� )�IYq�d�/��V��l�R�uJ_e����q�6I�����]�=Y3�j$0���Q9q4�tsnTc���3��?O��1g�k�{p��-{n�����`���y�����y�'6������U(  ������
����� ��V��  	N��h��4�G�U[.e4j:v�:�Uk�3���}���>j#cD-D%�q��\N8be��Sq����.���=����*m�����݉R�g����N��V�2^i���xL N�WtL�M�gCX�D_ hy �)�ĵp�J���j� /Z8<59��f���¢t\_�S?��'���%�-����Z 2
��jG7�waX_3�s���]iU
�ў1�
��ϛ����q�Į�f�%K%jV+���ˮ���7Z�Ay��[���(�V�|�#8{�O�O�uwT�5��=���DAE&)���Y?-�gk#0�YPJG���r|�N���Kj���{�ǳ��<ON硝�x ��O@��������ln�"�Z/덨�U˦y��uz�z�z/�l�͝�ǎ���<�Hk��zfŲ�����2�3n�ieq�}�t ��C/8��Ǌ��Xw�j���CZd�I���55�ԊQ��6���e��qܪ�W�O4x��AX�i�xm��F���vQ/� @j
�ć�Q�ZΓ6�spO��p�S��X�PS�<�P�#P>|G�?�1 b�1;��$!p��_�z�mW����N^���-���s�c�ev�u[�V-X�Q�J�jK���U�l����6^�z���N�d���8%ӨW�?������#���M�ɨ��9�J� �&-�����?�9�?���5��[&�:U&B0���⣨Y�1��)Z�`�B ��p���BH��o� ַ`c#gll쌝�?aC�#�6�JS5Ǝ�L�?U>�5����eQ�H�M��3�ȑXuax6��lt>ߩ&>�X��H�
Xm(ƀ(�ƈ�_Xn��f;P��G2!�d��A�uE����	��P�#A��ɠ%f��!�SA7q圏��kh�xo板au����;B��@Ӈ7��z��Kr�	Łkആ�x1�J?�B����ի�z�o������`==�Q���]��J۹�
�L:a�j�R�v[��޽Q�\M�jn@����I�әk8�H�'��"��d�b��6�<Z&�|�=�|�%��.�{wk�֙��/!p���:�VB<�ł���'��3)� 4�?_�����R? ��؉���@�Ɔ���G%_R�6;�7`߾��Z�����4�˗��ZםJ��Z �@,*%0�|h�Ӂ/K5R�m�iu>����ب	�H�Nw�l��ę�6���G�����P���gW�>�V�6�=t�J���S��r�</s�ld���Y x�Y�sg<%��.�v�۸/V � �Q��t��O"�_ Z����45p��9y��7�|��X#�s�e�u˥V��{�b�����*ik��U=���*��oo��J������׵�����r�7�H)�\���i�_�������6p���!�4���F�hB#�nr�'�جh�a�n����q��4K�-�"Sr��������8j�Ҙe3˥��]�;�w̱#����S�BUh�+����ΪY��C3BP >��je��8N�p I9V�ĮPs
AZ!��C�C�V��i��DA���y���ID*a ���E�*�F��(,������~;��k����s���������_/�!�}Ё!�F�^����?����ʃ�k�`~�����\��������f��A۵�J���͖JT�FD1�n�u��x�f͚g�]�j-�-��p��{�R�'��:�%I����)�p�7��LE�|&���[S>��(��S8|��帝��A�C�h�>��Xlbi~�z�@��V��^{Ķ��mլK�g��Jy������j%��LZ[{��}��~�)�4)V�I�'��B�Oʣ�������y~�a�TdC�Zn�y*�G �	7�+Q�l�i$����xEIp�q�M�Lo�O<t�4q<����&��$_ׄz�2�Г%#�E� �*�;��է`)�@�yF`p}��*Ĕ��0���r��B	��@l���.8|U�'������s4pﵜ[ӣ��o߶��ch�J8��Ixe�f�����M�Z�Y"�v�8U]��'�G=�{/�]ȘJ�z��T�P$T@��iGd����i�}��}�����00��(�	���&�\0	/c�jz�5e9��kG��d�h��h:m��wl�*�#F��$��g�R6{����B��J�l6��˩'ν0�������J�*��c�㈆�����w�C�1/p��7p� z�(+��8���y*#	���&�Fq�Y(Jl��⚊D�#Y��r$��g�A&6�|���0�H���r�9��W9�0�D������h��=�x��(r-j���h�{?�E�,���Y���,�oV+Y�2�Y�:,��rw��/V�\JX���L�ݪ��er9+�"���~~0j����z�S����d�˼`�[����jg4�O�O&_��f����K��f�vv���8<<��ZWW�'Zș'`�����W�� /i��AܫUy?-{��{�"�4j$$%��5��.�'��L�#3e�j�8Y%���w`���ݿO����
��^@4�v���4v� E,)��r%1�/JbGCb���K���`��wfgg��������~��eؙ!�/��s]{�Ιs��y��������4�dh:wx��܇���K��s��P����9�D���}�)��H֬\�bi�RP�UK��̯Y5V���M-�m��,;P�Z,i�x�^ۇ�<�\32���*cS�L���W��/t"4`��ɣ:�.0���
:=��9��������Z���}F��?�����2|�s %-%_{{���'�oނ��h�bkjn�b�`'QX�����>셖��Z��mJ#`�ʙ��D��~�]1�p�Q����G���?������Xv���ɘ�ke��b:�����%;|�۲y4#:=Ǽ�ϼ���/����E�PE�g}�$�h<<H A�?yF�=z���q��#f���>5/�]�	�36y�Xˤ(�V��Y�,f�B��?�.��f�B3���h���O����G��?~ꖺ�&�!�o~�o��@���������&3]rT���j����cC����Δ�o�׎>f�==~��Jf7π�?|.�?yʤ�x�?=t���f.$q�������
d�-[�£+H�bQ�z�=�ڹB*�&�v��qkۿ����7<2m=��"�H�!,��pp�*� �?8OTI�7}�fC^��}ʶkףv�s���ojL8�{נXʒ�&۹����v;q�ߒ�Fw`�@�3;������q��#N'���E��f�Q:�
N�@[I8�
���
�g���
�7=Ŀ�ᛈ�l����v�RkH�;|I��KY�T�ɓf؆�[��D�56��8�b��e�X���S��)E��:F�i��!AHTAx.o)�''>�/k�3?c�L��!������d>�
�B�f��zh�}��o�B`�ވ����G+�f͂������R{�e/{��$9�6V�y�R�d���8���9,�xZ���X��O</U��%�0d�ǆ�4.��i�z���ݹ���>dU��J��V��KZ:�b:���������[��٩�ٳ��O{J	�����U�S��M�ld���#����B��X�N��u��7aȹ�>Gg�4���RD���5�ym3���c�u�e&��S}�y�_d�
��)��i�4y��=4��t`8�u���J,@��<���=���(�¿r��J����`-#jzz�F���������>�;u*�&�yt�����G+�K:"Mq�^��^��ߴ�&
d嬘�z�*Ijjij�~!�7�_o�c�Y�q�;R�i��z7����&Fm_lJ�aB�9��C� 0�}�$�{��>��������:h��)��oHc�P,Y:�jm{=%ɋ����-��>8|�?R�/B���Ĵ��8�t�OC�ۢQ;Q�����}��Ϲa�7��S��$��F��ty���+�T�ui��5�wcV,e��u�57�؊U�,f��Oo(�G�m�稱��~��?��p�(@�ƴ'e����Om��Paޣ���D}g���%���T �����jժ-\�ȦO�i�M�J7xe�}m쓟�����Y�q�uV�>[�m�����Z�
�8aV������������y;�^{��?��J�R�FsC�]�b��^w����$�P7 T�=��s#D�j�rS㇘a�ˡ����|caRu2Z�-/|ڱJѱ���tٱcv�H��v����Z,D, ��=�e��+���T���s��
#�w`c)5D/����y�_�.~_a�}E��2Z��#�����xN��������>/�y�J+��M'�&mN-=�V��d�w�
eknj�dH�:d�!�1V���GA��د��Z��l��	����G��?�yg�r-��|[6��B~����:w����}���㌍�0�^��ټ�����Ŋ��=�ȣv��
�CB��.�?i��t�m�������xOo�ug��B�Rɸ���/�+.����Az觶{ד�L%,�ΈU���ռ�ґ�ݶh�{�^7�%J�I��ۭ�B곐�T�;������g�d|l��r�$��/@����U*v��k߷ݣH�u���{��6�CcOz�r���>Ϥ��(6>�����ƣ�Ȅ	�|N��Tq���F>/:8j	����C���b�97�g��v��\�_m�<`kW�g7���d�j�l��O�j�nt��n2��3C"��D@!��By�������
�l�r[�q��� ��@�6
UpaB&|���|�j�(��jκ�qő���sߙ�6;r䘭]���ѓ���n��K_��=��9�i_^�u���oV	�ل���}�-[z��
v�}w۬����T�:�a�R�q�%�iJ��;U�W��k��/>��� �$qू#� :,�Ph����8�}Ī)K�O5k�N򪞅b�'�466[[�A�����=A��@�ޣ�����o�z��$y1.�K'�W��;�E4u��te��2�yM�bcC�\�9{�e����h��%���=6X�9�ۜ�X��6oZm�*��kV+Vm��%6k�*+V�V.��Z����ӂ�G�� ���G�b�[�ƌku*�� �3�u!���T�_�?e?8�rΎ����`:;;,I+�xh��Y=|����g-�/����fϙg�x���;�5(���>g��m��zz�����[�O�<���G�q���������9z��zp����w[��#�y$kK��R��Z��7�<�4C�P��B��ҡ�����]��<l$6E�p��覧�l�z��b�͚�v�H������}��W,a�;�����S{��X���i��U��x�Ё�+_��]r�e~ppӺ񢋶�&�l���/�9�a��&�.=CY�r����-�0�c�S���+���˸�r.��Z~*�B�V�a-���/�t4F[y
��U����������*�Aa���>����4�Ud-���I�ɀ��i�pMeG�*(�.c>�x����E!ߌ�M~�9�����-ާ�E)K����՞Pb��
���p�O/���f�b۲e�U�}�L&,^1�>k��Y��*��b���:=s= ��Y苡�B�����2&���y[�]�W�������N$��O'?U��_�����'��&Nh�	�Z��=���Y�6Y6W��;;�RK�ɓ��v����rNM�O�3�x�VXt�G��,�}F�PՒE�?w�]�u���>�����]v�k=R���C����fX2��S������i��q�V������R�'�:��fs���OO������'�����r Y�7kH&,��Y�������;݁��4���uڽ�?d�\���Й����z���ꆍJF�a���osС�O6��m��^@G/V�OMz� ��9P��<(<T�) ��-0侀���h"m|���(�34�@ 
K5v�q+��ļh��V�ͅP�ƨ�`	�A�Q�ƭ�b͇~�<J H��Ґ?�s0^�c� ��:�� ��
�1N֌9�s\�N��t�%��4]���ֽ���u��C���D��*�%�,0"�O�흼���7sQ'���%��X��+ϳ͛WY��o���e?a��]��;y�����/��͵r������~��)g��⋼�<?
g�fCP��৒��g����}������ov�sm⤱�c�ϭR����l�v�9`k�����\���B�x�����=%S=j���Y���>���[���v��U��@�}�߰�/�`�X�����p���Y;r�U*��v�5L96:�ޮ�_�MMo>� @�����}׭��8��u UR*��%gt��J�����}����SGͪ��h0��X۳'8|��g.�����!�s�h(��h'����c��<c�={���;<�B~�֕$�ѺR�BQmz(�I��(xHs�ʀ��F#�� �� �!��Um 	"��Lt�+�O���{�nc0	��J{H *������q�"� �p��B�u��2~=�,�cM�^�F[����?�HT�%��c�\SV��������e�N8��p���u����+��P�!��6�X�p����o�8�4i>��x�ɚ�L�ISfz#u2���N�C��g7̅yt������-1�G��G�O�'���g�+�K�X��ڳ�q{��o�ʕ�l��V۽g��$��Rͪ��=���4���'\���
�U�yٮ={�'����G2Z��Po1X�{�����?�^�ɪ��>�����L}���'��[.�#]�A�G��ѡ��,"�J
�PP��8|��l43q�j���<b�o�`:~f�OX�T�LC4�x���i��費�}����&�T 5�3O�����P�\�4s���6���^�!�P9\�k�6����0c#���)o,�|G7�6�4h��@F�q�'j�*�,��QPR䖛�ޗ9lE*�vQ�d���
n����S��PU�b�    IDAT ƳH;}$@�΅��h.���q�
�|J�������o�;���X��yn�8lֆ=�ƪ����T9������2�%$������{�{G�uGC�����z�۴q��q$��|�X"�%�s��G�<�"�z�,I"g-D��kh��]]��=�Wu@��8;�[@YC�!H�f��e��٥p=����<��~������ĉ���m��KE�R��lޏ��w���2������A�����mFֽ��9��w�?�GkK����&O��η�n�S��Nul��D���T�:1`��d��/��^�җ:xP����o���'u����$�:����k�7��m�ڑ��<h����&;S��//��'�#��,�Y*�|$�D�G�9��I^ݧr�L�X�Z���9�3�|��_���_��_ٛ��&[�|���b��Ǒ��9��	~e/+�M�T4ę�( �
�J���h��p@�4K��z��4z(��c�gS�(W/*Jܺ@?��.!%zHt��*����BF 
�3o�>�����{�y�% ��2�����.�2�c�ŵ٫p�\KN%D͝Nn,��O ���Y@Q?E�ϴF<�z\h=�N�g��O�{�f�qo�N��WY<^�r)��=e�c��/k�c&��/~��*���O�;�D�P�+����i*���Y"�A��F�'��g��|,<�����8��}�~t�]6}�8ki�XGg�ˑ�PW(�~�C��ȱS���o/x���+�\j'Or���/|�N��v��|�V�YL�����&�P�xʶn��^|٥��sº�:�����8y�ʕ�%q+{S���c);~�{���&�_��5N�pҹ��ˁ���~���XhWl2{��A�_u���=Z��r6ƦM�BM��7<C$y��8j�	�$k�JIgw8�c�δ؎���;��;g�t�K��S�'1�#w�Ղ�O�UW]��� @���w���C{��"��j���E]��1����-��0�QJCܺ�n6���Ґ��^`!MYZ��q�9�w�;E��q�v���ʚ�`":F<u��$Ǯ��k���`�~Y%|�W�bQ;r���FAC�X��`3$��0c�,9��ή]�|��@�{I(���[ȱ�Ϩ7��G�,YC�LtMt]~
�7/��:�|:"��×f.O�}��_��Ų���CSC�J�|�y��Y������V/�\)ǩ�˜�7n�;~�~����zg�@߲�?�я:��<+����}h��h�����u���u�ú���l�+������	;��k:�X_o�^�����f�2v���; ��*hρ�(�݈v�I3���׿�Z�Ҿ:�ڮ�OZo�)KRʙ�o޹'i�J�j��󗬶+��!��D�s�{�8�}� ő�/��O��/��n��&w&�Y�!g�{��(�U����W�R�Y:�D2f�b�R�F+Wv�D���5wX[,f��p`f>��>h+��7�!lj����r�']�|�;��!��gy@���A�C[=r9(ꔅ	ˋM�5ѐY>��h�(�A���|>�;c D!�!�9�X�+g��|0���5U���" Y'����Su��S*Ғ�{��)J�uHj͹�"���s-�s͘��s4K5|ѳȂ���]�z���&\�R"��s��PEX���H�p]�IT����v(9o͙�>��Ng�)A��D��(E!���8�-K��J`�4E��.�8�O���~)�L��榘�C�D�O���|�i��U��(�@Ѵ�eZ\�O{�>��+���A�_��Я���(+KJ�g���I<���jլ���i���Y6G���G�Bɚ[-�/{��qc'��������;��A��3ٔf6jU�xh�H]Up��ۅm�9�j�����O~�#;��a�b�-�;ޖ/_a��l�Y�X_߀o��[�V�?8|�q�I����?���]w���x<l��f�\(���G�;�k���Y���T�fU��d��h?GtO�,��д"�$V%���U=�|F�d<�&Z?4����N>�ʳ~�S��tTϏ��\2� �Ќ �K@�"��B`��}��ph�'�y8�&�$� ,�.-|$��0�9��LBp��"hq���c�)��cf��G)cz��\�3�G �<��3���Ҁ&���V}���K^����p/��K#`"K.v�ʘ��ʕ+]��pD������sM9b�����d���5t$��{�;�\��9���5`mn|�y�����x������e�l�B���`�����݊�8|�	��˖0�Eђ���b�X�
Ţ+J�Z�&O�i˖��J~?�%�I���Wc#M[ʮ����u@�'�����W5n	tYV�=B��[�E��ﲥK���wn�n��~;~�;�)�BH�̙sl�ʵ^h2F��Z��o_��/��t��s��!0Z=6�Lu~�u��i�F����Bo�́�����k�X�&L�ds��3/�M$~,�& ��X���ȍh�lG�I�r/�o��o�q*�tp�}v=�����I�Y�R�)B��ԩ�=��V��_f��˂�l��V.#��8��WB	�fӽ�5�sڈ��9�����;�0ǯ�إ_��W�Y8�D(���@���>g�|�+�
 ӵk�:� ��CMH�A�O^UNB�+�xrσ%G����kD�5k�g��0gPvX)j�~�m�����6w��hx$��A�%�C�@C� \\��B����"��p=���q}� ��? ��e O(@+ׄ˿���z���گ9@�RB��<@�#��Bp���[n���F�+���A(�,W, ��A,� ��]����g��,��3��E���������}rMX#� ���`��=4[��ૈ�D�)�oO�2|G���[8o�-]�Ъ%:��=I���R�f3gͷ+.�;W�����)錒�X����=uʱ��y�E���u���/�gy�����\�
�8C	y�k_m��u��\(�Ѯ�v�P�𠱡�.\lc�O򂊍MM��?�/�v�ϕ�h�轢��^�4����$+��~P.��W��!�6��M�ߟ�����������?~Jq�lT6?}aqS1�
�\���_�ʠ�)� ��X`��\|z���_�O<hǺ�[KC�J���ͦ�Ix�۾}�=��G<f�B�C�jη���
����C����׿Ձ�g��׾fO<�sOhan���@q��!����t8�� _��v��)�2�4y@Q��p,�\��ܓ���'�=�y�s� ��.�`ܙ�\�w�֭x �	5B��9����T�y��b�/�uh0ƈ?��lXH 4���S L�}XX '�A���l�F�'���	��!8s�<#τpŢ �����ٯP��9����y�#�*G�o��o�}X։�@�s/�k�6�����,����1�&�N�}Ü�̿���ꂛy欈Fb��'�)����f�G��h��v4���Ϫ��m�ƕN��I_��j�wĬ�e��]�Ɋ%B&���|ɝ��7�C�;��n�[��H�?a�$Wz��ST${�3L�?���Žy�W��J�9a�Xߋ�Jy��Q(S��[=���;��g�5g=��h�6W������ji��0O��!�K���D�������^�>��x*�>��'o;w��~��v����2�i�p�ho�xh��o��MZ �D����}?�
��hh�̑���l���Б���Ү%KŃ�_���j���{~�����=�B E����B��ac��‿�s����::� P|ի^b�=�<�����h� 0g^8$r2����a����G ˈ�Vh�h��6 
��ÆF����%�!�   <րC��"Дo�sO�t@��v�o4~�eВ0P0��� P�V��r`�,��5f�h�h̀>ό���	B >�3�@�4N��5��'�)$F� ��AX"�����Cb1�>�����D�p},&����A�#�{"`���9�^��.�'����#9��� b�y&4c��Dp` h�OΎ"�$ ���;|)�P,���5K<cߪy���Z�a'�P�z���u[,�i�r��u'�' ����?�1����,�ٳ�z�7�6���|�c�R�ϣ\$@�yϿ�.ܼ��iTidM�p��v%�$Mŭ�ʺ�w&!pVW��b�����y�p�O��Or>�is�Nu�9cƌ�C���lX���~Sf�Y��ϡ��&����CE���� ���Pa��4��p�n�R�֒9oP�]���x� �}8�2��,^|�M�>���G��PB[�N���k|�2'X��O��2�(���������{ #a��|̫,$@����3�I��������Ƽ1���
���so��f
�:tȅ��ڱ�rJs]@���1���9�p#���c�q�C�kG���P"$������=� �'����~ m��S��Oh�B����F�h�PiD�(D���[).�`yp=��8q�<��ڡ�h�X8�)��E�@��B8 �/��s!�z���j��=Þ�o�`�Z@X#@x&�-
7)oӦΪG��9ڇ�ΔQ�$����R�Z��W5|l)��B��1c'�KVX2�h��R�Wt���op���|��.(YC����}���d�27��!�."���f���`��R����B��X����ΰ�E���Z<a}�Hk�^g5�_~�����j8�?�$�v�"M<�B!;�~����t�oEˤ��TZ��B��_��_��Dy��C��h�����-�q"z-�x����U=���Wky+�؞}O؉c�,ӀI�������j�,�ޤ�+$y-�3��V��h�?�q�$y�I�1 �}�� D��PCc( Q�Y/Om����������I����Y��]�Ce�2��e�?�C�p� �	x�
#�@c:s���4n@P�|O��1&��[�L�#��z ���@`��h��A	N\�ﲏ?ό Ch�>��2V���%��7�G��X�D�H��3
I�E� <PMF@]{T,4�dyvE�)Z�9�|ȷ�ȗ(��'�s�gB�����{�L�nY����O�����5��zl��e�y�*���Z�jD�4�،����ɳ����C����k�t���y�5��S�7��>*���<ɡ�{�_�A� �a>�'='ק�K�ۛ���!D���+,s�9E���r�����2���=|�]񩞞�7�nB����Oo4B:}����K[?8�нG���f�)'���q���9�8���X@1���5�{���G�R�Ǣ����s���ai	�fh��n��v��S������>ف��b�:�/�&R	����11^LN�����(h�������"��?h/4>Q��h��1�����%=��b�a��
	�o
)0E�ֈ��'�(��Xt��U�d�H�(�C�T+�� `|Ou\��>�Z��\GQR$����r=��M֤"�؛\K�+t�g��*���r�!���e�!D���h�|NJ��#d���?`�gEI��<p-��n���:��b%p�}��i����y����}�+�АIX!�m�/�u�.���_�ڤI��${*=�jP<��;�G��@�<ɋ�?
������8�U	���U���B��u���@���38���8��h>���i���@Q��4�)�&_{��f�������I�����fU̓<�0s��җP1����7eZ���wP�OA�
�xk4A8Mi8�������>��G>2�@h���*�v&��"a)KZ���L�b]'xI�b)�<���?l���'^�ڧR�;(�R��p�����p�vc����b>p�AO *  �Qx
��ϡBbJ����7�����[U�l\��aN�	3~Ɔ���@B���u|�4~w��+|
��;��X�@��*?@Bٰ��W������)M�����ݮ��{K8z_龾A_��q�����T��br�	�
G2t����N��!����G�Gs%��s�̫���{�4����SF5SM!Q�Q�$���[��8^`k�,�t�jTM�C���KmּU��W���d2�)-$t��hL{G0��sS��O����� e_�w�5�Y��`-�|� <j�� �J�=���u���zC�
�J���B)���z�s��f��m�>�����3j�5����^���
~BX.FA������]*�tS�8yN�IT�d� Lp�*(Հ���o�;~0U����UճZ���=Cq7�>5J0c2;z�ö?��� ��2����{?[�D�����/tǫk6�vc�\�y�X4�F�I|���s�� � Z<�,��CX��@ �
�s/zB�%��i�:P�'�4DJ�LS~���e�&d�E�1i_|A��4Ƭ���"��rUn�������wyN�/��Z�l��D�B��A�/E���" x�Q8���e �������J���a˜��+!-Ag���|f(x�<����tV��Z�B�������B��p���S$'g�-�իϳT�j�R�
��-\����_c�J�2���C�Fē�z��Ԩr>��W/G(Z=��,Z��!�'�H�#��u��ϧS��T=��s���)�����M'�<�s��030�'b�$n�
�w+�/�ԁ{+�U�6�{��O&��4�W��{�ő&�CqzA��E��u���ٗJƬ�����s�>q�k�P��H���G��w�o�Y��]F�9#��� �5�����s�n��R������C��� �04�Q���H?��<#��sv�P:�kp �� ��f�=_A��m�T���z)dt@��ӜųhW�\h[6�6����)U-�j�9�۬��󗢇�r���p,|����`�̠q�T�,�`�?���*��n��di5fBR�W�> i�I�=�B��C�����ʭ����y�p��B�	� n�bg����!rE�* ;!��<�B�������H&��c6 �?�hrI��a^����:���O�c�d/�J��il����=���
�PŇ����_d�f�䅹;r���ND�?��NJ]*�ϸ���,����m �_ڰ��у�\�g�5��'����/�n~6?�pc{��O�R��{�nظ�jeJ9Sч�кcl�����:ަL�a��YS�8/�\Ĳ��W�lx@������9T`�4{�9�S�Ƈ�#�NTD�<gIB9��"r�T>���Z
V�5����OX�<��?i�|��>;t.��s���?^�`�U}�tTN�`~�<��S�.y%P��K�e�e�G�;�F�Y��l�-( 'Ǐ�P�UG�v�P���u�I��Q�J՚[&؞������C=�	Vb68�PO|u�p$�!$��5�\��Q矿���0�I�����""H�h��Eل����^��p�b=Ȁ;�q�z4ƿ����* I^O�����C3�zd�mӆl�����ސ�X�HDƊ嘍i�`7]h�<�C��*UK%3�h@��$�|��A�od�K(��ɏ�)�Q���N)5�y�B('Ih!h!j$�ǕM|�жi�Џ�7p?K�$��J<���3A�NXA�w��\� ��0�j$�}���$�37�k#̐�I��Åz�����G�\���7�-V/�[�O�l��'��{�%�S�&.�g͘�tV�p�����f�����t�+��ꡉ8��w��ͳ@-��I�l���<�8;�� 9N�{�����ϥy*�?��C �vklHY6�m�V/���ά��(
"� �X��Ŋ�3Ѷ\x���!L
�'I^|	�-�s�\�5��;���9O�����ij�e��+��R*{���	-G4}�ߛ0�&�:�O�2�/����{�i��D�T��o�+�����'/� ~P���N�B�#a!� J�@��G�'`K4�����B�CT$o�    IDAT=��5f8��'Z�����UK���֫Ikk?b?r��z�I�}p�͟;��1�	�EG�F���ybŊP'��@<8B�������AU/�+��{.��sm��טkY�RZ��ϵg��2���O=,r����CU�T�,ޒ-^0Ӗ-_d��P�Y2��`
��?�2��l����b��/& V ���_��C�dE��E�I�Q��a��b�!(T%����G
������������ng�O=���n���:���$/xp�RK�)�Q��G�"qy)|���(� Z@��(���Ђ밍�Y)"M�Q/�ŦË�
��[�Zo�I/�L�(�&V�ZKZS�D��/x�z�@%[�p�͟7+d�B�h�K8y\�<�-�08^�|@�':ģ�Ik
��B�P�gb=���2fEJ�Sʌ�tT���2��8Nk�Q�9���:���Z�2��%S+�<d���P���Lc�%S���<�*U��:�� �zb� /�y��Y⥈,�a���5�.U��AqW����x(9%"���g���K0傥����O�4����G+�P����h�l�F��S�jH���-t�pnii�E�e��,�;�vR�66��uF�5��Q�o�j�x�I]���v's��}m�����>K��?Md���d�}y�1�'��Λ�%��//�k8�G\����o
܉���\����X1��p4ro����}�=���ϊ��"�c~Jy��U3�O�����>��t�Ϥ�V*g��9f-�)�2�+18�A��ĩ�f�z���cA�S�z
0τ�=�aťpVi�Hi��E�D�Jm(d�L��ǒ��CkS��\�ԦN�l���>Ι��<�4�87	���{��4N�R���U���b��v���`��fO�m��_�9�f�E���MJ��kRH������?�I�#�H�����iq��+��n�,�pm�6Q��?b��<i�l�e�^�ө�QJ�'v�c]����gΜn��~�3F�	��|.�WQp�����_q�K9���@��p��B�3�����g����w�OQi���?3�s>���:E�-=��Z���� �C5Oj����9k�]z鋽�o2I&P�p���!ڇr�p�(e仼���p�3�T�q�?����G��	�$'f��6�lkl�0���X�ʢ{���?�'�[���B�D����Io9+9��K:WC&/N�J(�If���+^�r�0n�s}D��S�N��\2�0Ƕo��}l	o��%�dh�
� ~�EI�UGvM�̹t���JV�^��b%۽�!��M�Ȃ��|�7N�f�ut���&%~��U��G (!e$�׭e�~&?E�Q|%J��Z��
@8ʔU���� ��Q2���
�hR
�>�@�E���~r�X�6�(��CNa�<��!�\���F����I�o9�d��}�C�+�\t"�a���C��d9�"HX#Y����"K�<������h�g.f�]�|*��퓴B�7�wX�ܬ��n+W,��X-�h�bŒ���[(a!�����;`�&ݟu���6Dӕ�^���W؟�ٟ�Y�B�zq~ɘ�ҭjT)L�(��m��\��Ək�=��'�0c%8�����;�)���`��fa+4t����Z����ꎢX�3M~�_do|�묥�1X�>|�v<��u>hM�F�=w��w��:e�KUK�3��J-6
�!P�v=un���S%�M�g�?��O�#�xp�>��{��ah_�x�v�z�N�8`�B֒�%c���IKc�x۳��{߃6�������i>2����hN!*~�vv�u�ɆV�3�B��E	I@ոK��(� �����åB����G�5%PD��k1&e�J�]	/�[��響�
�IX*ƛ��B�{�:�k�\OUe��7����s�R��e)Ei���sܛ�Y��ҳ�7����SB����5�	�_O��~�O��P�t*f�B�mް��o\a�b�ҙ8ͳ<ο/�9�Z[�ٺ�<ڇ��yXl,P���Tۇ�Y{���k�[�盽�P�-@(P��o��"�٦t���Y�\�\��k����<��,��#X�����^!V�>�
�P�`}O�'M�r�Y�u�֛�{z�=S���$��y\�)S�7_�*����V-Yϩ���#?�'�|�Nv���f���/�bp�]�l��^��#` �������
�S_���ԽA�!���fΞ�%��4
�C� 7R�'����	�9u�N�<l�~zc�V�X�XC�kk;����Bm�~(��}��3X��Z�lF6;σp �pg�R߈�a�J�^�q�?'�U�+����Ł�����Ɛud>)��f�9c�GF��!sH����q]擒J����z|���N�Q�D �_�� �}d���&L|�^�ʳ�ٽ�AV�E�����B�j��{��� �oX�� sĵm|Iܟ�9撹C9�w�&*/j�L�2�+�j�x�$.�mP�_�Ϟ�<�G�����S�e�r[�a�U����$�����i6a���I�@��垓!䓤O/R*�y�k��G)�����y6�d��A������#�@Nb)3�I���K����{�b��{m����s�c�굶v�&���%�Le�;��fh���BEÿ��ugga��[?���s�3|��aH� ݛ�'o|�l����kk�i?{�^���MQ�b�jI�!�j��_�%KWٺ���9����}����)�P�p��+��~͵oqI ��<hm�G���zmr�U�=�޶ݎ>�!��$2�&ۻ�34sɖ�ݤ�ϬuW����q �ď?��mkmE����u��9�S8(<֍�u@�������=���T����>�`��6�8�i��e� ~��O:�p㾔� �ɑ@s�z����cԴᙼ�s<X`���Yփ}��!�(W�㟱"����������C�s;�^MI���O>Z!�{�Y�ʝ�	z=pO�hQJ��_��"�3.������X�p�wXc�\��&h �%�����5#y��O-�b��3|�}⵼��x�fM-m���6v�T��˚�.�֡�C2c���,}~9��\������;n�Az#�����9�;��B��#���<��`A�R�q�i{�ч��'wG�1�K���z�5���V*�l` g���?��Q3�a�
��{����m���~8�w����Z�Z�7��Ͱj�h�>���������`��KK���w>W���S��_��lŮz�[h �]9�2���� ��y�k�>��O;� ro��M�D�i�=(���?Z��Uc�I&,�(Y���־o��j%�P��\��G���)�?!��_�X-�FJ��� 	��j��@?�Y^��KD��h�<� g�	 ����e��?��?�k|��?�/�@�i:z���ŢMQ�N�� ��V��F��É��`.Y�@G.�=�3`]L�:Ʌ%�)����\��hX.T'eLX>T[���vN�̯��9�K�y���?�k����;4|@��`�ױ�G��P�Mj!!d�/h@ ����{D�QdA�r�
?t"�E��BbL������g�UF�}���)�`���Z��֭_j����9#0n��l����a�Q!��]h��D�F1���:0f�����Vk<eͭ-���WzIg�?���X��a�{�ö�\>�O2Q�#��m�欄<u�{C�|��kv���,�����~�-Xx�o��|ͅ>��|RZ�(�svk���?� �i��ٟ�ɻ��a��}��ٺ˭Z�Z[�.���]��Y���v����f�tۖ���9|�2aY�K_[�G( 	��}�{���ń�۶�,@��06�\ФG�},n�Z�j�y��v�X��k{�
���
�����q����M� -6�G4?ټ<�f6���ƾ�-Fh�@�2ln9����̛@t��j)@{�'?�@e�5Lj5�ȸ/��T��µ��i<���+!r��E�s��d��C��-娱�кyV��5�y��_�6���ͅ@���u~��<��'w� �U����b>���p=,�xz#�Rv���c��+Wz�4�{
���PE�!X<(X!������e/1G졨������ь��?���D�V.[`�6,��J/x�����Y�-o�V��{�s��sJ�y=�9m'=������s~ޒ�}��wT�,`����+�	�|��{��߶���)T�N���o,�Z��}V*Ǭ�x��ʥ/�K.y��3����ӳ�i�r���=��붭���a8��DC�9m��p���J��:q�~��o��e�������ug��R�ӝ����l����6w�b�r��g��jY|�EW�q�U���e 0���"� �5����DȌ�Ex&E���:����y�
�~�E��D������i�_����
�D�'��.~_��&��w�.PD���`i^�3���IVh�h����g�xa#<�3 >��(�CA3Ѷ��];��� ���}����چ��h� ����}$˫\)�8xa�߸?��3X*_�Hx�G�((��K_�VԞ��#�lX(T<廔�� ��Iz%�	j@����}�.όe�����)8�y߳k��=#�g>��\ ���G�T�'�Wq��zU�P�'I!�ꀭ]u��߰�҉�F#��Y���u�H4[�d0�Xܳ� tѢ�&g�g~���>Ŋ͘5ӕ��v�g�Q|��P|�s��_؋�S�'��c?�x�-_��&�c;v�E%�$䥬�7k��t���v�D����`���w{%�#�N:%�s{h�?^��?��������y��m7�`�I۷�q��[_����V.�Yǁ=�M�S����Z��C��ڎ��KVx�T �k�Q���w%�GQ��b��C�븃D����>�P�3 "pJV�����Nkk{Ҋ�^knL{)j�留�}Z_��`i��l��YV�~$�a�W\?T�ҥ��8>����^��Q�]8oh4_�X>80�<��&�"(&N��3�	���C� � f��C �e_s�N��v��2� &����ϐ�?��$3��j�O�<���������G�:S��b]� о�7_��^1����h�?/�A�#��cg~^��K��_��S��茙�&X!(<B Z뭩�ѝ��
A�傰Ta����������B�Y�*���N^T�ݸn�mش�j��OTi��V��9K��������4y5\b�CE�������hwkݣ},a�}�����7��)^�q,a�S�	5��X~"�9�(��{����a�2�8q����J�Q�L�-�-��]m^|��'g=}y����ߚ[�Y.[��|�c�Ѿo���9��O/�r�Gz�{�:��_�7
Y8���Ʒ��g���v�7���������|X�j%i}�y��+���w���e���Fʣ��������B��h� #��Vv����v���@�T��/9w��y��;rp���V��Rλ6���X�ہC��{�L�LC�
Xϛ7'���k����+�ꪩ�%����'������n�Mp�j<�g����;��w�P���] ���,%4o�V�Z"�`'�1 ,C�i�p�{�X�y��o��8��>%�X#iϬ-�`�<�Ȝ�7Y�'�{X>�=����>��<3���������+��F�0G(���w�� �N��Rr��ޔ^{I���B�OE�9R�آԠr:Ȣ B(�i�U	��8�D���c�#fӽ�?�\���(���O���[�fm�ʅ�y�*K'jV,����V($��a���0�����uʜתa�]!����٩>4�P2� ~ᅛ}MX�T�jemI�"�G�����??w�z�~t�7lŊ�6}�T{��G�Z�'/h���,�h��G���d�'n�L�����ܳg��&���ׯC���_����~�<�d��Fx������w��55��Z�ٿ��?�E�-m�W����!y���~��~�ʵ�=^��.�
�L6a]8�?��X�K.��M4/�M��p-]��7����nΣQ@���Wԑ�{T�|�������U�$%��*W�6n�4{��6��COZ_o1����m��6w������r�у��P̊� j��U恟�gW��*��h�\W	[��G��F���j��\ �\��o�D%W)�_��Z����
��}�[���9�џ�R�38e�)7@m�J@SG�~݋uT8��y�3��5ŕG�A֏��T)�?��b�?p�T��	�g!c�9�H$���O�mUP�/�BC׋�c��14���H,,�:y͝��N^�5���Ջm��%��o����:M�ן�1�&��~�R���{��J=�'a1����[�p�Z�I�я~�[�2.|?(������s*kN������g��g����1}�577Z{�^��(��T�1{�g;-�i��ǻmݺ�쥿��Ǝ�d�v����S�N�?���[g/��F�`�1aM��r�6[�v��,���ʀuu:���]����J7ہ���y脝8U�����\�����)�8����H���щ���ܻ��ݩ*f�/��hn�t���Ås�}�N�Q��s�
�>76���L|�����x؎�pb��Ϝ19�i�*pÃ?�*�#�s���f-j`E3�=Z�Rq *��<)��M���P�: #Z/��?@(�s}����=s����氢a�!�=�/�&��X
<#���+ˁ{�ys}�+��s�;�Sy�ų�󀇚�3V�����%$��3�¼���{pO�Y;w˴�V�,��ʭ���7��2��J�����ESro������i�E�:�Z�(���~	����?w�i��U<�w��́���W,؆u���-k���'E���%l�l���j�/Xn�\Ś[�?�Y�����[��Af���!jg�	��Z��BAOr�yvĬ7c���p��+���'-��B1�:�3ꊱ�-�c��?o?��Þ�՛�����S��w�|F����l@��Q�&O��K�����N�b�8�P<ekW���\s�UJ9+���c�#��Ȟ�ŇO��	ո�eK�(���.X������㧲K�����+�� �N��p��׹�@4�����pM����f6���-�g�'��b�ϓ�0)S�9�{o�=�}��lt��l���6s�3JZ�� ��p�0Y�d�8q�/���9p�lv�`����������9<�CB� �t��	��3C����4Y�(������*x2��a�������<BN<�����rc\|�5b�rƁPC�#�/������@ �(�7~|!̓'dM��kϸ���S��d�TB�H�W�>�a~� "�D@/��f�j�0�`��٫Ap�7et�������b��,C	,��>�KSԂ��W�N��ГV++Hc~
��4�o��L��^[�`�-[���P�������y���<j�B��O�����ʁ��k���k�Tj;g��r�-!(�=�S�e��Q��3�l��U�}�־�������',CK�B?��ez��6o���n�fkjn�����˭_�g��%dߟ�Uo�r����+>������8O�f�KUZj�<���T�����~��ֶw�e�h	w�,�`��۰��;���,.�@4HT{��%��F� ��c��M�1݋E�� ��!���>�i؃A5���=�i�|����!b�b�s�X���V,�(ڢ��'���5�>h�42�q��
-��w�r�g(0E���n����K4Q4~g���l�� a�1�e�XHD�`#�=959��4s��7�a0�����D�0��:"��y;D��	��B���p����0v7B�8k��e�#܈���K4 �{�
 �m���5'��H/�V���A� ��׮Q!5��8h��J��u�Þ�E�;�'_�T��@;���ח��U��5foHj�D���	0G�}$��\��=b    IDATG�ߟ1mz��{���������T�p���^��S�*�����z�2��6~�Tki�h�}Yo�B�x�O����H�T��Q�z��#��"�e@ԗ(4YF(6��Z�`Ǐ�����ܹ�:vX:�r��YҦO�iny�-Z��b�����/~�KFU"�Fz���?ra7B�b�@��@s������:�?g�d{h�`'O��G:�6q�T�>m���0�
� �qڢՉ{�@�9d ����w~�@�8��� p�1�f��gpͬ}�>{�G�����U�9�N��Œ�u"g���x��*U"�ʶh��={�����5���c�U��o��Vki��I���p��Y �Z᪀. �Q�A��{r��	r� ��L��;L�� �ѦBݓfP"bEEf1���y��Qr��/͔�� >�q�L|r-7���C# ̱$�=������N4"< |�|��)��%�M��~��pX�V���yf��1��x��rҨ����s�8\W&�0峚	)-eq�Q�_�蜨�XV��Y~}G�CV\0�0	Y.<{��s�����P��7�v<Q���36ab�ūeKg���L�<O�P*ٔi���/���4��>�XҊ����T"��n�5��jj����'c�p�����|D��(�2��o�iӧXKK�u�:aǎ���9y��Ek���lμ��L|���;v�W��ekko�Ʀ��p����+F,�������F�m��������
[�t���9-^E����꤀S��O#Z�*5ʉ���&�Xt�.g`А(���녺�.p y��H��fO>��>��V�D�f2�Gi"���\���{к{�Pn�g�3g�͙=}��	��4���Bp�]]�|��PG�k�dx�MJ�����? bM �p��������NT��ׅ���a�p1.���4l~b����.f6�:V �6��pFx`�Y�ϸ� �p����j��u$�@���s*�-���`a<<'�\�
Q_�����-%�ː=��QA8��9a��o9��KQ�;�ы�����×����t~2�*�w&�"�)?�׿�w��`���'F�[J���p ���,
�u�{3f̪w�:s=��\�ٚU�m�U�<x��$Z��^7a�]��_�^M�c��A��),2�����@_���;�|=�?�>�x�;˺D��x֐u�|�+��+�!(����l��M[[�z�Fj��FX�߼�۱�I����G�p���)��;+�}Fn悃,t��@�ĭ��j�9k�4��.��6n\ocƵ���d/c��'�w�s�k�Q�5�Iy��k��B:|0�OM��W��8sB=���u}��V��;~f'�z;G��	�DXa2����~���!��@ uP��ϡ�H�l^�3P&���}�k_qpE�E��	��xf��d0��M����{�s���3��X U ��2P$� n~"��_���9��\��.L�Do0� >Z5c"��sPX ��'z�g����7�@p���\!w�5�8�@�E�>'���Rh����>� �b`��;�[�M�	��H/�.�0@��v�sF�xi�cBԌ�'��Ⱥ�x�τP�rGi��>e,������ʘk���sO���@��B���I{e(D�?�$�,
B�4iJ��^�?�N��n��ev�5���Z*�L"c�r��u]�w6v��Z��� F!�Y:�`U��jN�p^?����A��NJFdh��V2�{��nͣ,){P��]�K�㖑Q��]I?X1w~�N;x�@(��sX��b���j�Z�2i�gea���8R�#����K�ZM��%�Ny	 b�d?y�7���{,]o����,8��& ���������h��f`S����7Ra7�:�&>}�����FS���������?��T�
�!�J:��q�9G+��a'�u��� �E��3*MV5  ��\xm �a�E����y�&��� ���=�@�= D�����YE�p-�V��=s��m�{@�0���	���,kD�Q2�@�]����@P��C �yc�h�(? !��"���hrMb��h�0i�\��M"�9�惤D%�y< s�P&"�u�>\ۭ�tz����9o��~/�c����S�eNX�B�����J��ҳ�I � Z�5�%��q�?�f.���[�������X������R5�i+T����-8υ���i�BD�"�����7�)��66X���^����U��^�0?��^��b��;��Y�g��:8�<�´������Dw��U�EK%C2�sWü��[�ʒ����C<�)�t}ʋ��J)$	ł��� ��kj�;:,J:�	p���x�l���z�'k�U�������$�z̳�?��R��d����;R� ��4s�8
�s�eL�P���b�n�*iH�N �h��zդgNWϼ�.�Xڧ�4F��84�����gĽ2~Ơh �3�7��6�h�pW��r�	+��9S�-�仌��Sa��}$�枊����O8a,H����9�F)���h?��C�� �&;���yQq!���^e}��e���~��{�}�s/|-�e�K��B`" �h7o?�:%X��	+,�#�	�G`�Z`/Θ>�����!bi(��鞵5+��u�\9Jz�k"��է��isl���ij���B�l�J���S�롞��>p��Y���&R)+�r�V�/��5V������"��(b�>7D#y�!�h�4��M��j}\X�����b�����}����
fR�%;���j{��zCo���A
>��,H����^r�Ձ֏���D��P�#��'�[>4OBBh�7O�<�����{n��y��r�R�c���p��u�k���g�?��q��(ِ��IA���<��m��1f7��|q�q�r^lz�I�աW��(��p99��:5�L9�&����j��:�-�V��Ys>/�Ut
ϫ{i��$%����D"m�46�����N}nDo(�����XO��G�W���}�;4Hi�DXae<���^��1 HZXS�?�+�Nܓy��}�53��דlV ����ʇ`]��_���,�:8ЙX}�M��O�0Ux(�+����^�2�X�X�Z(�i�C�W�����ﭽ��~���v�4ѨkV)V��e�-Y��2c=��.^iώ�z
����	sa���ߛ��S��\�W�d͘/�rg:���9��N���+8X ^&\��H4�Z�{^<h>�P���(�;��=�L�� u͟�^�����Hl0�������F�_�%^��A��g8DD�l��B��Y" ������ 	������w���Y��S�*a��G��͜5���B�؀����w� /LH�=���V4:>�Ӕ�D�h�p�p4H9���B��h)�(� 0��VH"��eP&h�P9�Q�T��{P2h�h�P��JEà���g���c� Uċ(\?��c��l8kq�)����$��1C��S���U/��% �B@�F�Eĥ�S_��9�/�{(�ZV�@_�������#掝�����_[*�v|��I��E/r��ń��9��<?Bp0��r(i��ի9�%��4�	Ʌ�S�5�2��$�h0�/�!�G�k!�
-���Â?�/��Y.{�6mZn7� _��&�*��]a��-�l�l���Rҙ��U"D�Q�Y�����ł��
)4n�+�����S�J~]��{�H[]���[ �
_E�Rb����>�����3k��^v?��CæB�?U�L:���o�����$V]�ߞ���۝�� &�qSۣ��{��1���y
��Ъ�{�d�VJ�`:�����'�!�\
�Ā>�ihy2>��������"�	�c���w�#4X��8�8`|0g 	�K2���g�Q:T�D��!L��Ǣ"j&Q7X]|W���h� �N�(�%�b�B���1_�7@d�h��;�	�?�G\�U�q){��8]��'m�>J$����hd�?���_�h�]����O*�27�?J/�$��o��{q��g�x�R��pt{�{�A��G2�`f.��TL?���Ǉ�~�~.��%N^Ԣ�!/���b.�k(I���6uZ��sZ�W�o��C���/jum��/���J�d�r���/�CQ�������k�p����`�>)/�m��� {�hG�Z(��K�'�Gđ�9$1h�`�����?�_q����t��ax�B�Y��/
8/S�τ$�@w�0(��
�BY4`�)�C�Aw��������А��0�5F���@"̀��y܎�g�r�A�fko��K��J:W-4s��l4�_�9��V}�e��1���o�fO�����I�*��.��E2�J@��U�	`��4����@  ���P�8 �d Ѐ�*��|�*Aa5����c�!��.�
����3s-��  
�@�po��8H8�X/�<'U������/�3�����%? �$�ƺ#���!�g]�2UrӾ������lf�q
������Z.�����!�%��ĺ!�A+A%`�ܱ�]�/���|=��L����^w�y�3��ZN��
�cF0c�!DP0X;	��t����N���ok�.q�'Uݮ*��
��ҍ�_�zMj�s���רµ�C�p�cu��c%Z(�U��:�pܑ�߱�V��7f	�r��C�Qh(Q�N&�5pf�0Bԋ�&O��t�nݶ���==�?#�ӭǝ�1��s���>8xc!
Ӌ`�D�������%�@��()�;� ��h<����9|)���1^���v��n;y�Ò�rp�Vj�H5Y[�Q�羇O�%��?}����f�h�`0�n�r�cf^���ޅ  �s -<?`Kr?q ��7MH�͠�-��`B� ����E�>?4��5 }�w��� �.s!�8�l���z�j   �3r����h�|������R ��x&ƅ3ap	 �e H?����H��b P�)!�b2>r>��u����c8w����A���Љ��n!q}�A�s(�J��Y��,XM>������M����S�3{��W��khl�<ւ����{���G�����SXŬ#g��V��8�6p'�+��Wm�t"n�j�V�Z�߄�-��Y�Hᴄ5��n���Vs���Eע`����{0;��\{�gF���r�d[�l�$?��9�Bs�$�%�	qbSB���P\���$!�⊻-K��fT�h$M߳�>���=�myfd$�����5�=_���y�zֳ���փ���V�T�-TCX���gT�O��H �;FX���k��]r�O-�/"6 ���Q=����ܲ��==ݿ=2�G:��+�y�j���@�x$��[�lSo��2�'+�>�>��8m�U���ΟI0j�7V�C�vX{�~��=f��R*V),�Գ���n���������o�h1��gW��@ �D���-�' �{>t���j�i&�B��` �X�o�� ���%`�#��^2� �=��my6� ��� e (�}��z��K�P  ǳ�;W ���� ذL�2ѯciC}@��?1�U�eL� 	m�c�i�6�jG*.Yi���:�����^oL�PY�˟g�j�Pb��.�ω�	�b��b���al�� zyg,*�w������챋6m�׿�j_t�&j4�+��Ip�X�;�U�s��Ρ5��zO�w�����b�}y�x]��9��G4��iy��3��ʝ�Z֊�-\��.^�ROh�z�c�< ��w�>��	1�x�p`~�+��@��lO W�cx�����%@����޳����0'��6}�uw�z��O����G]S����+7o�FOo�F,d^��C���A��� �Z�c!1f�R�Z&I��t�^�SBQJ}���A"��5X ,e�q�'�`��g���^��XC�E*��G�7��]?��r��54R
~v��uf�
`F��k��ď>��SX� )�\�pŽ1��$��X�����R�@W���X�⻙����o �����Yx�G�`����c����B8�TAE<--tx,&PB����|���|��=��k��N:�X�B'�����bժt�(=��(2�O~	%��p�\�!��}��]�Prܧ,�����m�\ v����x2�#o��1�Yp��x�|�G��:V1��vIlǥ����546:��x���L��њc��1�v�{��Xg�#��! E�ܹ�O��}��O)f#��_�ފ�~�t:k�r��_J6n�$��%�Y�P���x���\�Q��$fG�/������|�j�:v�0j&�l�H��w��H-;�~Ľ��/`M�'#�y�hL����4�O	V����O`T�g��C�\(\�B!��{�sN�v�MwW,M�5��bV.Pf��_���f�^>/+¥m(��J�*H'~�c`�B[ <E/&wb�v�c((D��'�T��6s��`����G���~�|�q�>Fk"\I�y�Y���>:�x�G��������P��{Խ���s�9@u�X�܋��`�K������<;�����m$���`���^������ه�� &��]��K����]`aSo ��V����X�ܧ�`5����R}�����|�uJɽH�X|����"��y<�2�B��NUD��2:(+!�G&�;�
���/�Z���b��Y�y�P~|�u ̞��N�9�'xx%ހ��g�������ؑa͢������~g�w�9��g�s^΅7�K�ϙ�	�ּr�	ڧųy-V���,��kVZ"R�����K����[��l��(�� ��k�A2�����Ywoh�ٟ�YC*���?�Y����ƻ�~��+X�q��T�b����p9���?��;��1���>�Bry���UJ�S����ӯ���ۿq�Y���>f>��������I��Ix����CB
3�$��E��
�(Z�e�B���=�����h�W���p�'Mg�Jɚ���)cbx�-���v��[gW�����q�6f͜�Kny����Ț�Z�p]!X���y2���r?�G� �~��@�y"���z��"��ZM�	�D$�H�TJ4��$��p�s��¦������R�<�)�NV>����<₹GY{R�pn%�q/Ҷ�K��O%��̉�p���xMx)xP��TO���[��?��g��X��t�L�����c��b}:��#q�Jc�w}��>|/�������,�Jy5U�Z����� ����dB�(�J�8xW���+?���*��s�8~����=�W���6yJ��k�>��@\�x}���{m _�δP�d�¼L�k#�u����.������7_�ޗޫ�5׍���Ҽ����Պ��q��/���C"#�9*5�ϱ25�*~̐�w"?`���c��vr1eAk�c��p��sw=�t2�I�:���e"���y���
*k���$9�8MMf�����V���aY���:X̎v���V+��Y�Z�bs��O0y܄�6P(Z#�,zXT��/�ksg��C��h��`�t�LƯ�������
P��1 ���Ƶ�>���'H�*�zЕ�㗼)q٢K4Yd-�2Q� xn���6r���i��z�N�,�kl�V�����{l+jMV��1����_sl�A��������D�������Ρ�J\ �
�'����*��#N�	����,f���pn-bl/���#!�/�E�k�Vc;t�X��˟�2�C�"���7׌5;�F<K��<*�w$�oȦ-_豄ap�,����2����%2Y�4�;����N�����U+�iCRk��ݻ���@��\�x�I    IDATt�E��>��Ϻ�#��K��]=�%.�-�m��ܠQ�o���E_�~P���m�q0���ij�X$�6�yG�Dj�k�{�m�Y���}"0�e�9h��e˫��=�iC�,/�� ����yйm�|� ���-�1x .Y��r�ha�� ���@�i�X����n--��ˤ=��#.Q��g�Z����{i2�I�d���ϛm"Ji$��m���+� ��T)�p<Y��U!�wՕ��U�&�����_]� �_�qh����\T���������-eYr�L��D5Z��S�|��k�z�K+s/J���U���[�eK֠�x- <S��v�8�<C DupD;r-��� d@��>X������N��I8�Ȇ�������u�ߺ�)���ϖ�П���w�x�AV���<h3f�t�b-��L-Z\;�t�p��"������}�!�����G�8O�:#J��,��v�U=�.�i+V,0�-���܍��GgL�n���ם�)�B��x���/�r���h����-�_�ީ�o��g�3�����_≃��/hl8��lC:�S��J��?z����$>��9�*������?�Ο`�T�o �믻��]�B��\���bu�o�ץvP��;d�q�A�z��]�jչN��8TO�>��q��yˮY��Cf�iY�X������c�w?�%����)ƶ��_J.D�aGfB*8�X�ҭ;���{����e�>D��,]�O&e-^�ʗ�{�uC UqY�ҀkR`�����5�-��N �`. �w�EO�k$�C�9��L.��J�d�s<b$��4��c��*�>x����y(%���Ȋ��X����5h�g�q�d�s\���E��hav�2R��χ*��Q򉡼�
��=���r���=���s�<�V�ȸN&��HB��3����1u�+��s���i�?�i�S�Ѕ��r��p�5�x.	���)�0<��S�k���Vڅ�s��{�� �$V�Ž�������K�a�W�������@<�"���&��1�������[�t�0����cbC����pA����d���t���93��<���E�u�ڈqv׏dw��c���b2u�4��?��$y�V�b���NϘ6�9t&���|�2���O����x89
�o-Ł���y�L�@��Ǫ"�&:���@B��A���B�`;w�ԺzY�B����>�����ms���^�9�o�J��}O��W,d��:�Fp�[Z��D:��2�wJ2 �h�YXP��FÄF�$���Ft饗xP���}��>� n0�8X$ @*Or,�E�)E���J�.��a2�h��"�Ċ�o�&19�2��*��;�����-�<=p������Ce�M��Y9/|0E�xތ��	 �x�я�t5Ǉ.Q|����F &c�w�@8cL���`�h��x�=��� �\Ƕ���R�s�����B��9��do ˟�� 7Ή��kg_��k"������c�?��յ"ϲ~���=�l�?b�;рıh�T_ۇX��z�{m��e��5���v�o��J5n�R�Ə�l6n�r%�u~��{�0�w�g`���_��7���j�f�t�����"��2��x�4|g?1��1����@��qD:s���y��<[�>�e2$�%����=_��sx�!X>f��N���@�	N�>���o��V�<�]�|�߶m�x�>;���z��2$-�M�.����3s�"SU|6���4�L8L\H2 ���f�Q�< �Ԯ^�[��b�wv�ֶ�V��F�5_�5��%�wo�=��v��F��h���7o�!۱�h��y���C\�	�\'���@� 90�lQ��< ���H��&�{��# �dâ�\,,,"�+��)��YЋcb9�|Ѣ�3�X�XX)�`Cͱ� �(^H b�}�+Ã�<o
�2Ӹ~����ɽ��&.��<�7����ޟ㑸�+ә�)S ೨�����=� �����G��F���2�E3��L���ճc�O��O�y>��V ���?���?���YE�?��sƻ�9S��g�"I5 �3�(����wd� ���q����T<ԓ��k���˸`Fyĵ����YWح�����X�V����;$�H�$%�B�����l��ɶp�
Kgm0_v#�󧼇u���4��9d/O�1������w�B�\�2.	N���sc�+��{���x�믶���pgg{�=�����S[���7j����k���um��3�Z�y�����{DQ����=}u�[F��|�)�b�6n<�^�ZR�y�kn�k=|���U����)���Ҩ;oG���ŗ\��\}���I��Z�b�P���L�s�� �﬉	0a%���j�hR��ԋU,?pܞ����
��Ɇ�Ka��UϿb�X�-�P��U�f�(�P��)H��|Os��

���ʱԙ�ߋ�@����ŁkYu�yVX�,�,xz������aq� K��,(���� ��U�p�u�Pٖ�3�Ylx)�6,8�EZ��]�=ۯ
	���\�!����,"\ 1�����0tV4�b��d	�+d�+נ��|�'��C]���b
Xq� sWO�{9�a�0f9.ϗ�Xt� �� c��v|xWlG�>j�o�y�8�Œ�(�8k.Ԃ%p�ߙW�'ȳH�����1�����_��������v�R۰�����K��l��6}�|�0~���|C�8/��s�_԰�+���}��N����*6y��B�x~����R���7�)��*��n��6��?j��6n|���Z��>5{�寰Y3�z����vo'�{S<��8�7����nX�����k^s���a�%beoܞ�Ĭ����=�2J�R
���{��y��b®������L,'��QCrԣ�k_�]@-�D �Ky��'�?n�Z��F&`��e��n���\*����=d�����w0wsm���,(�H��������d�2��` hi���bun�`u�`�tx�,�,?��9�� �����>@V�,,HJG�i`U1��o��(րE�D0��(�@k��%p?瞻�3}ѕ�;�Z���k`q���Y�w}V�g�ǀ��҅��?���y�O�p�Tw�= ��
� �Kޢ���G��R*	L�N�g$�'�<��}d]C�K��s���ȣ�X�޹>���'�%ZJq����}�x(|`����y�#.�{Q@�,�������3�k#�>��_���y���J��n՘M�:�V�y�������c晐��F!�9i�|Ǽ��_}��LG��l�Θ�)p/�:�Zq<��^���&����֪��m�Σ���v�Z;�d���Eڑ�.+C2��|�M�8�b�?����n��.=WŉN��>�7s!����N9���=�o�tܲ��v��mͪ������u;ׇ
������:�TN���.���_�T8@�)`	������2�\l,?TG�v�$��W� �Wy��
�Ճ�J�j�׬��նm}�ʕ�gf���}�?��J����"/��?�#����\3Vu6��4�@������p\,y����m��� :�29��������"l <�?�����e�1�U�sJX� @̢�����n�kp��_q����{-N�3�[���11���\/ �W�g�f%� �b��xlâ(�7V?�f��9.�ͳe��&2��3U��.�lx7�[ �Y����<S��8d9��c9��J��$�,2�I-��s�/�c�O%τg�"ʹ�r@�f�xx�.��=��5��X$��)��:��Q���@
,�ݜ����;Pw���\�qKe�֬Yj/8�b������N�l���h�:+�Vȗ���?���{Tq4zG�I�P�ǎw�_�t��� �����^�;�`Jf��k�^�f�C��'�s��J���wYC֬�1c��^�� �:�I۵��i;x�î��[v��K,�����[n��C��zE`=tZ����C��>Κ1����m�R�;c����.�� Q�:��A����~;x��
Ť=^��3�z�D& /k_*^
r9^:�@%K +x��+\Ѡ@�`�:`r�^Փ��[��X��a{wo�d*XU�.����'�)���ޖrΜ�/��~��w�&^�g���w�4LN�^Ԅ�f�� � 7 �}�Sn�����-]�@��W2S�K9�&�hY�R�̤��z?��z�����-����{��e��j{ (1N��Иj��9�ԓ�e;%[j�^χ�=�
���?��8���zO����;������ ���H;B����kd_�)T(q � �Y�J��}���x��w�޾�6]|��Gx'�>X<�b�|����g5����jW4u;�x{Jv`1�	P&��P���%s��;)�����Jm�V�^b�?�;y�����'m���6k�Y�m�b�A�Ū'|�H���Z����j�x�c7�ڇ�>u�L����s��0�0Jx&�R��ϒD�K:l����lŊy6u�$�����BE�*I�q����=��6�i�����u����.>p�e��[ Nk�߼e�{z�Ӏ�1d=ׂ�ꬕ+�k�bM�������wϝ�i]�r�==]��SM�u��:b�r�����.r��������I�t�r*2��v�%�A��h��i"^�R��v�x̺��z	
� Z����t6z�Vk�h�"�3w�s��:��_)� ���I�A�,T~�"����lϳ�X!�: ��.e@*�\���\+�	@5����� �&%?9�~��nط~A�5�'p�3Wb��Zt�VO���X�ܯ��h��4.��K�(J�d�k�X
 �3���g�������pmx-����XR���Y�Q9�!��>ʑP�-4���1c��9'@�5J��R@����� 8cZ���?~�����&��H��Ϙ,
����h���N^��_��=p�,��VZ2�j_�z<&N�yα	�g: �C.	��D��D�% �?�2	�֗��dhlø#���Ž��c�|b���!����c�����b^��ҙ��ݷ��w�_*F�J���iu�����U��� %�@�홝;�ٌd�������_���~$�'��@]�t���~�*�A��;f���U���-�(��C�^��C��y���Z�Z���g����6zEJ&�� "V�^:?���I�$���䤙|���0A�(�������jǏ���������K��V�V2�4��t$�t�Yͻ�-��_��{*��k�v�zB�Aq���J��W� ��7�&)��ǩ�(IJܴ&���kW�W�e(p�'V1ϟg+�M��.���7ā�� �R�7�=��^ �u ���s~�'���iw}����u���&�/%�AaQ�=q��C��/���
���g�;��' U�`�B�Op�hX\�<���Pw,4,.3����q-HCG��Y���P2caN��;���KGa{��?���\7�� ��{�_�����i��Ӟ�5`��.�u�V���Z0�bi7q�e'Z63��.\l�Dƻy�H��:�hL��;��En��a����~���Q��������;O�4����-����]v׿��F&����{�b��Z�P���n���$;�v��{�?�J$�r@/�ݿo��3#����~�-'��t��9:�G2���'؟��y-�L&fw��5[��L����4�Vн�VM[_o�Z[�Y_�:��v���}5g��+c!��y�v���p�X����#L�%˖�%Ǥ����'���k��y�+���[��m��K�,c��7j�qaSm��N���G��)� �Zd���hI^Rp=^_<�:�Q�A�l .�τUr��tU?���J}kC�� 3�����A0y�K �v��n���@&zH�E.�ߎ��f{BD��[y&m�L���ST	���y�,�sX d��3����8�8}QW�^-,</>���#cDIO�PP�= ��P=�G�t�{#hK��uk�V�<<��<c/}��\����ze��3�ga�������o�UW��v ��?ng�\��@_�_������PG���3�S�$ׅ���_F�F����?j�dS1/�p����a��V)S�'��3$<��Kem\�D�p�ž ���&"����X�c4��'<N��/�ߺ��.@`� �g<d�~%��%:`�C�}�uw���i�N��q	g�}��/=a[��D�юu�lٲ���o|�Wm?��ϲ�H�s�� <�
�}N[��rOo�5#Y���2Y������k�s���-�(Y>�c�����e���LZ{�1k9�a���]�~�Ox&�*�r� �,� V��) ų���z�5��f"�J�+`�`%ԫ}F��#͖��,�1��u��ke�;����;N��e��/=|�J��fd�g��A�@8��]���� `���}q,I�ا�W��z�XT�J7��?E��L$a���(��}�p���H��[uQ�e-(|�8�hyql�~,`��⟵���!�h��`�����t�1��la�S��\��L��3Bm�3c�I1r�w<L�	),V+�`qs�LxD��.q�ߑ�@����}<+%)�W"�}��@��(����9�#��|���'�u�E��	�s�:?Q\1WD�`(��G�?���p��IXn��6n<�.8��}.�z&�]��U�)ˤ�s�Eό�{�^껇�����n�����qp�����]>G%&��ȳ��"�Q���=r��j%o�>m���HV����/b�4%-kv�h�5h��#���׽��]�֟ŝw��^�H�^������vǭw|����O��F������s�J{ӛ�h�j�*ł5��}{wz5O:��=�#��r�j=}�6}�"������PP�0�Eo����pR��A��2q�wדg��T\B$�N�T����	���
Sg春�p�Tm+�O&	�M�&[��#�u�;ޝ�Z?��f۲���*.$����җ�4��s/Ǿ��<���Tő��JR\���x,I,�ƢW�5��Q������U�< �X�Pyj�V��%/�-���5�/����i.spc,�47��.�l�_5� @Q5���m��F=D�`�J�����򈤢��&�a�g������έ��/����L��e��\���[s�7;�Y:��{��)��Z>_��	�-��X��={f�{�Y����<��cV�e0���e/}�{4ܣbP,N�w�������� 7�Z)X��xd�7EJ��
0x�i��K���k�T�]v�+���,���v�w=&�4~¨/�����?r'/+�X(���dMM��7�ٖ-[�u�a\�~j�g�>x��ʅA�t�B[�f�-;k�uu��D�7+�8I��ݨ�8���bB�
���:�k��+�í�:��y+7e���C��eqf�@Y@��i���5�B�xͥq����Ŋ:�c����_�Q Ɓ�J�~�,}��Jn+M��U}(Qr�)�p����+�l o��@ � B����j��n��nbN@�a�@7�v�;�AX�쫚F�2�M&�
}���L�;�ʊ����y*���o4�w�'��b1gMM	ה�� �{2���Ǜ9e�91h�Z�-j�`�s���Q��8S��jN�U����_��1<}�J��ŋ�Y�R���G�g�v��<J�'����Xn��]`��&o���Νv�Wi�EU��˿蜧5�o޲��{z^?���A���6A�3��3,��Oˁ����a�r��Qyoά�6k�\+US�8n�[Gdh�ؖ�@���ѷ�V  9'.9|,�����p��s�d+�7���ܼ���v��ak���L�EI�1c��+�c�e]�F!������ٳ�����\�,�_h���A���׌Sh@�PG0� l� �
Œ�Øb�3�P����L�|���Ǌ���)!��Ʊ��}�    IDATd��3( ��İ��U<�le<���ù�sa��	��"�˜!&�, �$u�D�wά���'(�V��8�}K&ʖL�l07�q�b��U�����d�r��ͯ�T��K(P��A8j��"������e����K�͛�h.�u���dA�3���빱p2�7����	�m��&��hs�Tow���y��p�*X �v�-c���_[{�W
�Li�<�Nk�r˕�����G��w�R��8m���nx�M�2q��T:�rp��8�b�W�����\+_�=q���FH~�}�IU>���KC�OQ����/�=��ּo��ckjL�@H)GFa�={ۮ����������,���&U����_�q�}d�364���+ �$hȮ`3c��R9 '���n�ɍ�N5�H������C����!@����>�+�CX��`�X�ϖ)ٹc���5�qCG�m)���I1?�@)fS�aQ]R�)����Ϝc�z����n��B�l���v��K�j�ު�bE =��gΘo���׽�s,Ny��d= �M�
�>G�����R�7_�V{٥���"o�k�:QAAeW�9�]_�}Ӧ��W��M�8ޚ��=������;�=��*�g���]{��-u���V��
ӧN{�i��9�埈k�I�Ʉ���7a�xzQ ŭ��D1Şsv׏�vK�~�,�X����[IxA�̠Ɗ���2�ؼp�1b��8J=�������ÛTSԍ��Ɔ�[X(V����~�����4�F�������w�������w4�7�lKD��ĪG#KRk�)����θ����PQ&v>jdþ,���>�O���� ���9�Z��k�W�q��^T�T�q��it�*����?�w�aI��
A�#`��QI�[�ϭ�Op7?�kk�[a�6��Ze�j�UJ9$<V��l��i�f���ן��x<.J>S��8�;��٧����3����߱��\ڍ����9F!:h6���ޕ��w������gKsY�	�%�Ugj�������:ފ2�k:ʍ��QhdS"�ͩ��
Or���x�R_�\�[xJ�����U���^�X�r5>�w��f����/�8~�%Q��!����~ ������]��Ԑ�d����Z�&O�a�w�;|���2^�%Ȃ��NYc���Ͽܽђ>@A� �C)�\X��we3��A��Po��Fߗ��#� f�U�o�Cy�Mݤ'�x������Ko�tz�H����]��M�<GEtǠ�%	I��E��C�t�2�z{{���O�
�# [Dȣ1�؎E�Le��� z5s)נG�����e�ןe]x��}������U�I+�)�7��n��-��>b��������K6��9-����ɖ-Y�^W�ҌA�*����爸$��y���z����&M��m���m���~�۾��t����à���{�0u���{�m_;y��:�o����a$ڇ��In�/���χ��^ld��ł�=n|hP�T��g���g�a�A��EF�/^8ٗL&0A3,;t�X|(%+�a8�?�붣GZWW��u
�T������.����>cV,T��3�r��NA�i��>�\�G���� ��3�c��&"��J�%H�$ aٓ�Ż���[(E�( zz����F���L#C���F���#m���,]�؟8���N����u���f��Xx�7d�/@!�9�^��zw�(ܛ��p���}�h�o���]�ܥ�I�?m˥�%��mʴ�6q�6u�l�x�Ű��U$�<W��p���_�B腲m�t�]w�[\�D�B�c��k����T]&)��d�޸=HxQ��B��,޾�^����8NC6����YG����X�V�O�>��;n���s>�=��ӨŇ�������+��O |�{h���Ui��cM�	�y�*�'����PJo{��<Y�	"����8zsg���K.۳w�l�ci��5ҵ+f�-�v���@�!��4v\R��5*�h�_,<�r��{V� �]C4���
P5R�0�@�` ���ᝳ?��{d�����V6��ˌ���Q�A�@]Я�r~���&su���A���m����!����9�z�=�}Y����#*U�^ݓ��|�袋�f.Á���s�]bm\�%�)�H�V:3�.>צ͜�u�JU�� �Hy"�'yEy,T�$�듟��Z���0���?�C�Kt��xv�R�@��˳�=`4��;������a1�ܳʐC�])�ĩa2\v�� ����Sq�/h�8��Fo�`�EE�"-���x�dM2y���O�#� ��=Ǻ��Ο	�d���YC*i�b�R�=vؚ�m��`�/T��7�������T,A�o-�nՓ�<��>�k��Ac�?i#�O�7��L����"D% �ÄfxY t�P<:�<	�m۷{�0�' ��l��>ۏ�}��ӄĵ��2����#���k�������V�^�F���G�g�>x&j��v2���`�?��J����͘�6��[��x�b���[��9w��SU/���x�Y�h�Z˗0�2f���d
'���)�h�nN�,��������k|��dqkjhp��8��uq�м,�F.�� 	��àO,h��GH<�>p�ӦO�����O���WC��?XQ-���>'�?�(E��cM��S�f@��M�H&��Vw&21QV0iFj�k)�,�IXS6fmͶw�V���9H`iii����r���' �MM������g�M�集
�R�@���ˇ�i�9��rI�b%3��� Q5O7�zD��*�xa�3V��?��%xw�I ��A�'��A��5r}���#g?U����b"��}@k@y��T
פ�o5�q��lq��^؍���f�zB���yk����˽��}@ۅ�δ�γB9$m�jP>)W�d���[�fNd}ui�O}�Ӯ�w=?%�*�ސ���l�G��u�<���,D;ɲ�1�^�e�{{z^7��_�h�jH��S��:�w���y�b��X`\`�9$e�äQ���n=�:&�Aޚ��{��J���"���J:?d���	�f.�梪 �<F���������󢪍� &F����82��� b��f���j�˂�*�e�Ŋ�q��1�����R�c��/-���5��kb��9�x
[�|�&F%�|��O�Խ����	>��I�+���E^F
s��(~W�!�9s��U�<�Ua�lM�[�֮4��:�SΘm˖o�L���-Rޝ���ۆ���%T,��{�ֶC�ٿ�,��bL<�P�d���r�(F#�&>G��O�8�� j!;�9Nw��;==��}a�����q��G-�ݯ�h�l3a�S���	,��ކ��U��D�z{�[_�u��Xww��#��-��v/�ݢf.���cD��⎁����5۠�/���2���]��ϻ5�A�hJy���Ϙ�8.��sw^���<	�r\��0�j����� {�(�r-c[Mdؗ�p�x'�cK�/V=�\��U�f?ߑ�����:ߋ#�~� �[��o�?��:Q��|�]x�9v���Z����x����>c�M�6߲��4N�B������s*����v��_}�
Q������K�+�K�bj�=*3S/�74���TOp��_��� �#�8,	ύ��~�Gp�Qd�);W�
c�KcA�Ť�����H=�X�i���f/�L[8�QjU�L������9m���#�왡�`T�v����?a�_=�cq׃?�E@I!ۡ��~�; %�q�ō���
Ń��lT�)���u�b1��(v���B�*�5J^T/�"�����!�W�R�;*�W)��Iu�D ��y~G�I��\�ߓ���������S6��a�
۰�\�T,���Ӻ�h�����V�m�}��P%���뱱Z�z�����?�s/��s�e$*�������Y��Kp��8��:y[���~M<�8#��u��~�7��O�	����?/��	�	��9y��M�ădo��*����:�8dmx�#}be��4:�V+)��l2d����0�Z��]���W�VP��?�\/]�����ON]�z�5M=�C숚0d�:hᡂX�
�dT�w��'?�I��_UQ�i�"�KZJ-@��2b|J�L�d�q��|Ϣ��,>��1�@U�gScP��XD���Ăǵ��S�d��x�������[����U+��mݚ��s��a"Q��W�	/�R��m℩v�K^扑P?(�<W���Я�q���J*��� ����<s� )|FYw=#�-C���Q^G0>��"8�;n����Qi��_��
�ؓ���xl����Rɪ�U ��B�8��� `��j��J�L��R��j%�V󖌺a�g2m�f�����l�R1���^�(8c���	�����>�B��,jh�C��G=�g\�DH��Ģ3�yM�9s�G?��� ��t��\��e؇r�xxT�e�����g�{�g(���8 ���F�-�	E�ꇅd0�?$v�����im����4�q��\gϜ�
�� �TUO���&V��m͹Km��gӧ�ɚ�g0���\��,Y��ZjF 8����[���|�;߶� �er����Ӟ�v�~G�GGY'�.�8��<�>����0����N�~�wo���O�濽���|�K�Ї(�@������Z[�ڑ�W���;��L��R�y�ZD���D3Ed�{�1 ?g�֘IX�4�HH�'R���ޢ=��6�Xƕ�R�-Yl�����Β�����&�#g�� /T6/�.�'W.�A�( ��Ή:��/2QJ%3�<}j�6���>�5��h��泟�ĳ�	�B���'@�<�*����8@�)>`�J��liJ?s�|��͟��,Z�9ǎ���-Y��ҍ��:	�C� ��c�P�͚��s��k ��j�����p�;k��P�V��,�t.��۝v�����~D��'��'���=P���l��[-z��x��>�/��)��܋�BA�u��[&��� �L����+7o�VOo���|�V��54f,ח�j�&��uM'3�
��i��fuB�����ِXLLJE��sTkE��+�<U*T��x�6����'��9f���V)�)`Ԝ�,W�)�,NF �A-n�.��s�vq�S|���:$9Tp���r�)J�׬d�_Mh�տ* F�H� �s��l���7Nd)��T^	�C�|�!���`��}��c�(���7��M�|�9�dYTH.���Ch�hu�W��NU攬��J��C�������?�����"+�������k�xUO,�Pճ��[�f?@���V)3��r������M�5T��S�[n��ٌ?��ɤ�ko�굽h����\�/u��� ���}�S���� ��5G<_.xŀr��� �΢LǼ��;�rȪU����`(I�ChH3�紶�GO�%��j^��R �d<e�]�R�;g͚��D�]R���b����� <���pl���冻����RkA&�5���C=�t"�T��;����l�\o�%1KE�Y��L���~���4�f�'l޼C5R�����I^����=�3������>��Ɉ�x�_}��սB%�i��JU�D*�ႊ/Z�e��y�O<���a�w��.6 Q�3���M�8��А�_)�d�B}�������F�-�xy�{�;$��PB� ��Y.�Г�8�k�
�˸Vj�qȠ`,O�:���s��	���P#��ڄ	Y;c�xKF�J�B��b%���[`/{��f�z�X
��q&�F����t� ���T&��	�x0ڔנX�EmK�Y�P�!es�Rq�l;�앎3fd�!���7`;w����l6m�R��r}��~#Nk�r˖Q���p��usή����y����'O����ϼ�C�����(����i���z�������D��FI^���5�k$��'|�l{vo��{�ZB�M9����T�|f�>{��m��M㖬��;g�-Z�0���b$����M�uY�xp��p�yNyB��ū�>/�	8������s��P�����ࣨDIe���ܵ���n鲅������;�UvA9c�����[�h$,S�%X�x��G>2T �kW�k;�:�Cc�{Q�,�(��w��]�HhA#>k�[�p~���퓌�N^_Tm��œ%[y�"[�z�{�rɒ� �4aǘ�4i�m��+㖈g��o2jd�blE��찏�|�{|�����k��z1�H
ʜ��G4\}�r	.��R���mΜ�^��Z-{��kjj
yh>X`����8�U(���T9*�=� ;����ͷ�t��i$�-jw'�Y*�����W��[:2�r��^%�h�;����O%A�ep�t�'�����A4iy�������+eȜ�J�����^�:.���������'��6�f� )��2��Fk9p���!���[&KY�͝7�� �.X5�s����������n�C�!X��5�d��A^4��;�6���+�:E����=`-�d���J��������c���a�(XI�h��D�W�,U;�Ia�����իz?�C�� �9�K,W΁�c:�V�7d�3�Pq>-Ķ��\%OX�Tϟ�>sf���z��r��֯[i]�֬�w�'�(�X� 64N��7\��o��P�Y�3��vx��ԧl0?���^L���8�X�'`�G4�(-l��+^��v�K/�d�R,dq����~2�T��=r=�rr���1=��\!gY�Y��?�W]��+��=o1�KE��)o�r��+�寸�z��z��c�;���O?��4M���sV���o�q&{���R��LQ;��XT
�s�Ԁ?�1Oaokuݶt�X������;P��С�ֲ�U���(nc�ۻ�m��O*M ��<���#p	�U���e�SٝJ�g0�z+d�X$FRA��x�3�:�S@ �PGG��h�W�,��� ��w��k��G=�K��:(�DUZ�	�sϪxn��f� :�?��O|���:������+�Я���b�@f���y�{���.��8 j%Ā?qU�9�S���D'�@�b��X�{�!����q[��L۸q�����W=�Z�ĬTIZ���I����.�rm?}|�ޛt�-�,�RZ�����+(m����K/���Z���ډͰp1Wd$�w��K.��z�o���J���ჶ{�km=d{����x�2[�t�-X�ĦN�IPK�����py���S���:�����v$�'��I��5kV�u׾��zl\cʛ��w��F�L��'��JO�\�
%���앶x�
�\H�ԜEY�L`$Ȑ���CC�[n�ś8��-o�^��eM`�SO��H�hW��9ܺϊ�ǭ����./�J5���mv���Ya��/���m��%6�l�Jb	��4�*p�:!����� rq喳���LX���G������f<�A�99�+��h
�!��{��?�f{G�, 	��$� x�y��\�V����Զ'}�R���BQ3$�\=��0d��/@H	
��P�;�g[>�}�˸b�q}����%m6c���|O�H�J%)��kk׮���W�%9+�l�3�-�Lv��3M6c�\,Z�`p,�^�i� ?���t�v�H{�;���hx)\���h��s�])�':�wB<d��q��gv��n��ͪEK7d�!��\>����	S�׮x�M�1�E���Wo��:;)�w*˿Z�>u���e���-�����s�H�IC��7�卶t�|ˤ��Ҽ�J圵j���nO��S"��.Y��{,W0L�;���>�$�Pޕ�����?��ݪbB�!�]�U|��x�r&&ނ,�z����h\�l"c�Z�b�۳o�:�-I]F�������m0t�( �9�C��e���^|-
�LLx\]^
�62��    IDAT)�~>��[^��ƌ�� 2H=�(� {���3^X��,7�|�?T,�_� cE�)�鱦q���0��Sr�cqn�	 �o.�.�?��<lG2�T;�6~�lG�K�$rn	*�RK��@�cɰ��Nr��^�YI^!˶��$��D���3g�V-�������Oٔ)Sfۜ�l��Y�;��К��\�`�����B���s}��G}�p�Ϛ��$Ç8���L(�{���X�R��Zﳖ�v����k�X�\�*�:��*��3`�J�~�^ms��̦bw|�{���ĩ��-�jq��iם�U=7o�bOo����}�M�b���7ؔIM�L���߿��\��K&:�<�-&D���6�׬�Xɮ���p�&����ʇ����qH�-��ʾ��/����E�B&�it�gܬ�kZ��l�� ]@��a���Y�<��Fk����1���@��X"fK�-�ӧX�B�PO|4�_*�MLZx]�E�� �	��k��?@C*�1�O �!���W�@�<C!z������\<���, �&���/�=���|q(��3��L�c����;��qh
�V�����".�^J5z�b���s}�A�ߡ��XCn�)����e��"2v$�4�<�-�)���騼�WC�
���r�f�2���s�F"d<��Y��L���<��-_��E�]���"�z�s�>������&���?q�,��' ��w�.��?�q��p�)X���m{�^K���>|�r�3 ���í�֟+��`ͮ��7m�y-��؃?}�n���!I�H#,j�~����+����{ð�O8�lz�2{���n�b�Y�h�����K.���B�k��:�&����m�uX�����}�h�
w�x�j��B3��Q3������2���Y|�!��1X̸��h� ���Qy�ᥞqK[��ʃ�M��%����`��R�X��w�p-��%K��i��Z�I$#�?��kf�cyj1�u� �[Dfn��H��ol��'��d|1f	��H.[� ��6xdu��c�d�m��$��.ՖȌe���� �l��N W	d=�U`��9����A�qY8(E���������op�d�K3Ͻ{eT�_����F��T�_�تs�؅���E�Vڂ%묯��|��QD�0�jV3J��	ć�|������
���44��ʜ��	p�k,d�Y ����v���k������w�[�l���h�-���<{��W�kw���nhN�6׮�������<������7�w�g%*p�G�X-��,^do���J9gG:�O���]t�:ˤc�ܼϺ����N5Z{{��,�h{���k/p���!���Sn!/��c1`v����,g^��s	(U��p�O%_��q)�{l_�6;ұכ��h41n���y���	�Ƭ\�[�Ry��5�KU�$����j-�&$�- �1��/n�I���ǳTޅ��#�@��ի�k �xW�?���G��]%�i!����'�!�?5�1t�E�w�=�`_��j��,V|ǘ��e�3 #���^ƍ(%�˼`�S������v;��ɤV)����K��ɂ�x3h�E��;�S*�J�l�������
R�[�\�_�xc �Z������#�g��'/�6�������@E<)��]��kw���v��sl�����������;h;w�l�dk=|�*��}�C��K|�o>c{�����ؕ�Y��)U.����J�~;��a��/�`/\g�B�;��	L��%����n���m��|�*��UW�}�{ߐBCV>3�f�r�X8X>߾�;���HT�� ���p2��|�FI�����юfk��g��#8U.��4Xs�ѡ�/��ր�,/ i�W��(	�[t~BC�09�������H#�?������L� `�2� fx}������E���w˾�U�vޥ�����{}�R�����'s��{?��@/�P �ԩ��`,b�
�]�{M!�
Y4���!�,����ˁNT�<��Py�(���o"^�b��֭;�6]��9�|+����ON�e�W�5�ĳKZ*�`�\�
v�P���'>����V�<ө7����@"��C���K�Ƶ1���b�o�������s�^lS�N����T��d!_��{Z�\IX�^�TR�я��������ܼ�KL(��>��l�o'��e�L�2�>��?�Rq�R���v�7l��U�y��փ^���?�tο����Ÿ�i9f�6]����kM@V�5�U7���7�n��@D�`yPPj��[Ա�57?cm���ԓ�.�(Y�"�Z$i;p��ԓ ����A�|*�'�%Ǌ��U@˟=E#���(����� �����qw>���ƫ�3�/e��r�ԱFh@���>���fl�p�, +`��z����?� �j�����[�@
G��)����˳y��}�f�6@kB�
�#��sqN5p�����4~J�gSc�����V�E�y�ԓ��J-m�M��i�d;���V(�,fiK$�<���ϸR�8������7W������%�Ur��ϝE<�tv���?�|�\k�fl���n8�����\�v��o�x֎w،Y���kǛ���:p��-��8O�����n��m�}���߾�ە�7���皑�>h�����h�_�-�?�j��=��}6�����`_xў�D���l9h�����]w]�����C�#���G��d��gR�s&�{��׹��-�?,(	8�H%���쩧���foW�M'���Ja��	z�v���<hǻ����=���z��8��8QG��:	�"Їw*�s#�`� :�Dy��~���=	EX�H/���*�ޱ�6�S d��R��&���]���O�'�:��O7.���E��wj5�1X$X��s P�]��(s���i�GM�J%cV��_{�'yŬ`U�7$wR�N��K_a�Z��unt�X��ڇ�\�Go��3qy.h x��_�5b)�7�����~N��G�w�0�bǺ�Q[T`qj=�i�]��~���k�`�7\�E�ܺ;��o<'�o�A�?}��n���[N?��r������e$��lX���]�Mv�k_k}�]� h�mmV*Z&s�����~/�0q����W�����V(E���o�;n6�~Ǫ�A�U�� �.#:a���z���E��re����b��sO!1e����b�<��-*b&̛� ��%�p�r�#���)��U����*E��$Y�����g�i8�
t�/�MI� �(�>@�"�o��+I^�Y$��*����0N����2FQ��v�w��E���)�E����N�`'�㆘eh<�c>@��!p^<%��1^��s�Z�	w,Q���Zb�֞c�t�*ł%��n��9e�6s�W�T+�ư�Qǅ�8���˾���9�so�L�ʰ�s�����S�#۰�bPʥ�#v��>��hsj���R%����H5X�T�;�Y2�`�����S�{ىo~�[�ӟ>4��)�v�������t�y$�@�/�\qk捿�z�3w�M�`--{m�Χ�ۭ��{(U�K�Y�m�s-�j�����N��Kd3 x�b�o�8��������@F�dU+<�QGh�^v�*�56em|R��%"���$���Y�N��Q�ki�|2|�zEQ�ꑤ��3��=�p����τ�?��Á?�*�1h��-����1E���0��'��z�� ٗE�W�I��%����3�n���߹�[N�`�(X,%��������@[��)��?�#��8��L���;�4*�2�K
�z;�9�ς���ȅ�&Mj��&{UO/�Xt*��05����T&�4Y���c�]In0���Ɛ����3���:���-���	�f���Rgh\6iG:Z�8���;�����^8C=�����%�^fM�B������/���	���- ���mw�z�WO?���>^ځ�?��^�y筱�_�?��?���zmǎ�]�s��O��d�̚� �R̃��H��%��ÝE����o}k��?�4z����?��?��L&ܠ�����?\�77�k��X�T�$��(Z��)�ʖ�d�>�%�F�^������j�Q����_��M�ZU%�>
62�Ƥ�?������v�n�±������^x?P����{
��E� +@�g�ƍC�d��J`c1�P�*���n���;h#�9 �𦼁<Z����������Ϙq��ba9C�2W 9�sB�: |����I%�CU�t*���>������:}W�%~=.�%K�yrd� �<�RԎ�gt��a��_�eμپ�>��%ܻ!��c�!ཽ���y�HZD=zĽ�'�|��Cpl�˯Y���=w�M�8œL)�����ǝ���t=aQ�$�1�$M
�8���T�/�d��f�&M�	��Z|����n��
�H�����>ॺ8r��ċb03�xXE�_�YX�d��
ϯ���`��m�3��b��~�R����
�Wl�S;�)�b��*D�����$��(�� I�	񏴃�B��`5�� {��6��O@�Z@Ř�l����h�js9o�5�v�\�9- �D�
�R��*�'ޞ�]��Ї>�/Zs>��Cm�c<��p�,
@ �x��P�?�$I�i�H�/c
��j$�
�k�܇J���Ϟ17�}�'qkkk?��1i��?g�$[�p�UJ�fR�P�͛�{����W���L�T�L���.X�Qt-�W�5&Bc�8��x2�B���/�`	�=�1O$��MQ���\�%j<�����$�
100�`WO�3�|X�K���7�s������-�e3Pqu	� {�ej��w:�,2q,fl+��Fݐ��=�)4�*U���X;z&��%����ޡV�];�c��<�Db
@R�/�g�a{��^���>��͎���9O����
p���ͽ��[�'���;T5��0��?���ͻ'Y D��0�G<3���w��|�� 8�� ˛y�1�'��Up�xrP�Gq<��}�W��@P���W�wE�n��ÜQ�"2��:��Mg@s�>G�mBL�RW�y8��k|�6h�Zf�_mF�R�X"��$ǁ���k�lm�Ԭ��B	�Z��嚢��2��_�����Qo�y}��/�o�>扏0���
/H
 ����3\��c`NJA�*�2Hهg�������JMwZ���-������Ƒ�J<�1Ȕ.���dnP&/������->�^kؓ��2�M�'��ŢW�� �%�TUO��F����3+ێg���P*��Y&��~�P���Q/�Lc5���._�$<Y��OF���k��^|X���\7�/W&E�d���y��7������ċ�nx��HOJ�y���&y%t%�_�+�|��R���U�Y'=� 0���1��X�(�THF��J�
Us�1$�Bu�6� |�L�W*��E�%�W}!�����چ,�����β��g�b>��wN���Ujq7�[{�7�
�@������y<^�Q,:<G����s���<&�8���Y��>�яz��W�A�<+B<8�����3��𼠿XP�����d�c�?
F�
�UISJ)%���jG��s*���ZH���AY�|��h�نA�W@�Z�u�	��*�'��Xaox���4�8ٵ;ةZWW���{z:��U:��������w�O�y��b��-^��fϙZ�UF���LV=i�%'T"�\�z�y��' �V�, ȭϺ�������"eч��pT�$8q (G@� c%�L>�ˈ#0�⃪�0��4�G���ƈ
�i�H&�W�.�"���o|�ϋ�EP`9]ŠU��/�|^�W�7��%�CUφlҊyJ�������Z]�>V1yz�O�4�Θ:�/^:y�)�q��>$-66f=��2����н��w�*j')9��j� �澸O����IU�ERυg� .�=F�:��^��H
���P��JӧN��4�z���K@%i#��˲R�h���|��>�C��,��n��i!�K�Ë��L�b�xSVw4�cB�`�H�y���\*�-V+Z__�<�ú�[-�E�@�Ѥ:�e?��a��H����-�g�fOwz(^K�j�s��X5xUp��&`�*�� դ?�e��A����eA,�n�
���$�D�;�� ���Bg����{�2/�`̊Ҕg��\΍�1������,M
����;D���3��x%|8��Ca�V�N^�U=U�٬X����t�rܪ��%bY�5�L�4y�54��L��
%4��~PBC�[Ro<ݛo�Kf�ӷ��Z�0i�'�a���H���ûG����_�Ǭ���L���^f��,m%~1�����j����������#�<|�i�Ղ ��� �@�`��~y���$��!@�Ń�G�n3����眀?n#�q��[�qo�ސa ����Xs�6��h������;CU�\�b� ��ϵ9s�[ie���*�~Z�4�����;��k��P>����C�/�%�幊g,�D����AF��V�!N����ƽ��Z�%ٔU�1D����ǖ�,�EsPF�"���b�x6m�<T�M�ζ
rj���=Q��,OEU=CI��4%ɻ��ϱ��?Ǫ����9�;g�^`����Tz�W�-�V$^���{�*������O9��
������|�	�X�h�U�n�h;C�.�AϙsS�D���/�N����2�O��W���)e��B�W�/\�.^�"��Lhd�������Y˒���-�4�xMx=h�D��;����IKO�[oO������>�S��w����'��b�x谵t�"�3w�U������g�
xVr�5����+��|�O�J>�
���>��{��� HW?��g��ƶ ���q���b�y����U�K��~
��#/�G�D�Z�W�2�D%�k�˜k����Hj29�P=�J)�}NJ:��a���a�ٖL�Ӄ�l�|�*�:s���d�s����H� ��<����3_[�a���}th�s}����
��QZ�1�Ƚ@�To�K�g�g�©F:||���UKގ�������M�z���?EwM���������{��]������ٚm)�R�Bh�iIDEE@D=��S�v��;˝�������"-	M@J	%=�������g~����g��eg7!	p�/^����Oy��y+
/?��4[nHic�nt]j'��Uf5��aM�N9�\@�� w:@l:!k������+�d ��;�c��L˺\�@��ƣ�-EG�Yˮ���?bd�U��D��W�o_��&��q�1P���������\9�����K��AZ�\RH��z�=�G�,;eq�:��\~<֛�#���La�tMi�^���w5�rƿ�y��|7��9�����!˘�ƌ0m�1���H��4Ǝ��c&��D7�`"���L���η.>�hU��c���+ĭ@�����r�����%4�����+��!���z�o�Ĺ���_�O�s���b��kim�����g��_B����
�� �ߵ�\ʙ�d�b^K�T�F͞��c0}���$0��Lw�:y�N��G � `qa�{'�/�+��ͨ�9�#�X�~��e�ǳV"�g=��7n����n��O�lZ/|~�����C7�+��G?F�<�2�Hu�J�R��7o�|��	�.��8q���-��;����m�ē��r���g2�T�Z:t��7�+�c왑6b7�Dp��(�,����� �����u�x���0�F` ��4-2���T�沎���5��w�)�OO���D���`�UW]�g��>����زy�ݻ�ݽ����Ne՘�葿Z'�@0
zy�Aq�V�Z�Jf,��9��Q8ɿ*��/�3�F�Ў����-��M�g�-r�PUgvЏ�3��S1�e:1c���1�D!��.�E�4"V݈��&6�    IDAT1�(+���l�p<��+s�y��i޹RKU����,k��x����R.������P�/5p|�n�zj����+-_�kZ���埓�HDҚ��f��ڠ�!��Kn�~�ݐÆ���m�J�}�D
ȧ�uTU7`��Mx��g���ΰ-]�ʍ�EC)9����R|>��[�v�]mh^��څ�
_��&Rq�T'`nݺ�������E6݁3'�S���O��"/�;}A�
Q�3E44�⤙���u�+M)�ƸX���mZ&�=͖^�[ɋ  *|����O�'�F�P<D��4�!�/�2�����|�L�S����ez	��wU�������_T�qoLA�C��XA��Cy�K�����|%kS�2	���g�ƭV�L��9�I�X�v�Pd�����ӳ�z����,�s�F�P�@߱#?�k�a��V����g��������i��=���'��O�fl�(0��3��"��aX�p+�"
�(3�`+��n$q1K��\�$�:ȏ�y�6V��4o5�SXB` �oni�~p��/���3jk-2oZ�I�B���r��l�
�޹�<_ח�Gn%	 Å�@/K�)������?�ً�h !���2�Y�C����6nي'�z��$Ba���p���1f�XdҎ(�ii,ء�G�
��:}h��v�Џi15*�����ػ7n�?ӧ��I��ǍǉӧXrD8��c*r��,�ٜz��5��+����c�f(ȇ�A��`v����H�6��x ^/^�{����'YR:KTV�>PПn�A����+e�w�V~6.,C�)3%�W1
�L4��*�#)�;p,3RE;��s"{��2�'p�e�_�p�u1�U��#�w��|���j$��رk7�T�Y�R`�Xv�:
�T�hXiL9��<��޹ۇt]lh�c�W?"!Ge�HvPkl���k�oτ@����$��#hjn@.������ѳ�s驝�Rɜ�|(���'];Ѩ#g����`��b?^��!JQ���tv5D�Λ�"W���4�
#p�e����"/i�^
N��i���J[J`e��xj�fJ��o���6y�
�tM�k�tHiJ�R���S)~��?)����N&��N�F�
WYos[�� �H!V"���#hjj���G�豣1��s0bD�-b�&�@G�������7~S`�����%1O�����r�e�oP>eA^��ٜ�1�Ҏn�����|��cu�ً�Q�8sYa[�q�- ���:
� � >�w�gT����}O�K�\b	�D��*{/�����`���x�����N��[
W&�᭭8��3��:�t��+-�i`X6L��u$n�D�P��ތ!	����{L�����a@�]]��gFO�˸ TU$�t�?\L)�"4o�SE:����k�{fΘn)r
R�`��,Z���v�!��"+��O��%�,K�x�����%ȿX阞�;R;��[�>�j��x�K�;�t�"38x��딿�wޏ�+��5��3��Vz�W_w��������RN��}l��4����Ǿ�ml�Ej�|�|i*Ϣާ�x�/���ۘ��|�����t��c<s{�g]�[��7��,�h�z�����wߋb!`����(��DCat'2�j����t�"�[�]��j�c����k��I�����5�� 8��;X<��q���G	���~N����>��!�����b�ݟE^�-�7J��܋L�t�����(䄾�k0m�q�1P�3��}o�ހM^���b-�T������|ģ��r�x}��e�9���(��ln���<�1�&q%���D����5�*�����{����ꫯ�s�������h-��4���f@2�s�������o,J>�6��������]>�t��b3�ѕ��3N�[=�'uD >��7(��u1h�̸#D�~��]3o~`�!��?l�� P(&m3�Ǎ&R1����#9ʡ�;��H#�A��n���Q�,��:�*<O�ŏb!_ dϗ�q���E����X�
pj����ek��Ϗ"��C�_4�y�	���2W�sW���S���Q��A�g��@��5*�2�.�r��vr�}�qN�
�f��h7?n�
șu����}d��d���B
���(�Jb�I
�5k��?]��_˥oz��t_ݟ�{��ʲeϛO���G��$`�u���<�����������u�7p�N�gL���^ U��woL�g��{Nq���8��_@??c�n��P���TWע;���K�3�i�%@K��>AG���5҃��?��������\����p���"��D0����²�F�le�y���	3����)S1|�([l�,�]�|�M
?�{��Pr����j��U%�O~�S��\ ��4P���'ٙ
*�i[���Ի`D~CUHrQ�r���]XR��~_+�+R+�
sA�cˋ�H&�6�Q�E�y f.8���,V/P0.j�N���Q��[��aaN��l��,'��;>��ʆ7��;>�}j����̆�.Y�
l6��X�h�)�%���6z(2�iS�dQ���&P��p�B��}���s��2�>���RiLl1�$`��������i��tPd!R>ւ�|V��/WcB���B1�N�0���=8ͱ�w���~nŜ�)�.�bP���kɕ�ci�X<���_����w�{�:��c	jn�l�*d�7��dZ5}Y�
���W�p̵_��A�We�]����u�x`*~׻�X���	��.{o(&�z ��^���fR���O௩�K9���w���a��عk��SScƏ���3N�~�������sK���O������:�ނy?��;n���,���8G�>��C���LC۲e�|�Q�;���0�����ο�ǉ3Nø�l�R@��G?*7s (35졇�x��i_�U>w�\9�L�,�O�� %�kA{ϯ�a5�8��6H�Ks����ٳվ��B*܆�a����5��!g-n �Ԇ��#	
�S{$�dm�>ט��:�l|SH r��M;��A;߹-r(�]@�.��.�Ի��&
�a�%����	rL�%�����/?r)���!�r-q|d�p,,�C?p0�xe
E
K�E�\|��ˢ�,�Hԏ|��K�_��~��s`��Y9� >Q�	U~���06W�sI:�Ɓ�E&�:�����
~�r�oB�ד
�s~ow������(���|�w�C�	�r-վ�/A!�GkQ�@�W�C��*��Ԟ�P9u�)Fa�����Q�����2�g�����g���n��I�Mwa붍xq�2�]�Y�c-��s�4kƑG���M�X]$���7��'�3}5��_0�����gZ��ITǪp���ٳ�J'��Վ�;6a�ڕ�XҜ%v����ޑDC����ך�g����g�d�YH3�.!���z �+'����ȇ��\���'��``��kj�Vֿ�x���M��9��,�ȣ������hf&����ȕ���g�,ɥ$�1A��1wF �l΁-�P0Rr�el3�	v��c	�sHf҈	�A��	������cڤ ��|�H0T�hx�Q d�����~ݿ$t|�����YՏ*ӈ�'��I�܉hU�	��6|���m�Fb�:��Y��C�e`�-����y}Z]�R�!��v���>��6�����|_�o�~:>G՜-�.����.}���o�G�����/o~(ʆ�xȚ���ۓ��������X�E�l
��*g�����4˂+Q�H����)�bj-���B��/�Ӂ��ͣ���ǐ�¢���g>��F�F��R5Y)Oz�����>S>?���5e>�B.G���ذn��چ*r�\&�5��b���v�L�s�F�Θ�/�+��)=Ͼ���1�����ߏw�o���S�rݼj����$��a4�U�ww�S��d"���6��&����۶�D2�Î])\r�[q�Ygوs�٨�����G$p���[���Z;"�Y ��w���hCie�@�/ ��UN����t����H�ՍƦZD��X~n�u����[�)u�+~�3��O],�@Е�s��s�s��;���Q����(Z��I'�� �pO�����\�֚�F��Ӊd"��a���]�W@�#Lh�K&��8] 4�0���sYz�z���6�;�C�lٺ�R[Z�͔D?���_&ldb<���	�g*�A$\���v�wU�0������%�3�``n!]
9���v���)�ڣ��khmѰ�P������u���;�mn5���F��b$�j�N���o��xI(Ïp��d�w�Ecc���e�0Ǎ�fKZ?���\�,�0v��_ l���xD�Ae%E)�Rp�n�Z?X�_�Ϸ��(��8��5Z4	>7��I'��/����g?kV�R��\<��<r�n��ғ�2��y�F��1���-�͛v"ѝFWg�]~f�<�((�)��寑+d�)B�m�q�n�_�����U_!h��Q�F�s�������v�0��S���ֶ��7�`��lټ�`5V�ۍ�Ǟ��~��f����]�(���G>�[lq�zR(�˿��� >����~��D*gn\o��P�}�9�����|s�<'�e�П�!�u>��[�@�B۷�㩿����{pͻ�j�'���R�r�_je��H����K�੿>�a��8��3Q[C��TbOp)�-L�n����~[6n�I�gb��1�{b_�B���{�X��R˪�d�YhF��T9�aAD����]���>�V��g�Css#�:�4C�
`�8�A:�3Mه4�LWdp�
�x��'�Pi⤣q���/cq(���A��OR� �q[ :;�x�'�Λ;��KY#ΏO!@߹��KMxؐ���������SO��L���5wV�*��P���}x~�Kv��SN��)cM ��a�@�IQ�_)S.��aǮ��랽����X<����8��	���o���;z?,����5F�C���s}�k_���>����Y�ϦM<�^����FMT��ɿ�c�D;���?b��ᨭ�F�Ƶ���0���JᕗW!k@[�5v>�w��^�;v첖�[�mvsPR�z5��_0�{������E��TL8f<>����V�Z�g��N<a��v�؆T�u��ՙD[�&���qL�|<>������I���B!S&ӹ����'�P0����C�Z���Be���J�/]��WҾ��M�.-���@��-"�9�~��Im�\6��/��IG �ڃb.m�j_>l�`A�b�B�y�`;vv��G�!���/��p��@�im�&�F�`�|h2S���kVo�#�=�au�p�[/E>w�}�8�R>f�d���?��#X���q��:�(�3=�{�=��.��L*��}��q\�΋P]4�`UU�4g��JUz�e_۷����?��#G��K�"_ �e-�)�r�&�g9dr��b@�����59n��v�t$��P`��#닙h08ZL�62�B��r���9gOGsK����Dssn�S*��*I>G�y�V�}ϟp�)'cƌL1��ǥ�z}�.5�M!�!��%�-�O<�3�:S���v H� A?_�b*�|ϴ��c��v,Z�8�	��yfS#�Z\����^% � �� +����-1� �����d	�%��#F��v�l��n^��L����-Ƨ����OE��?kּ�'�N�6MMðr�ˮ��AgWk�lB&�N|�����_Cu���.������+ʬ�ڻ�̟!���>Ǖ}��q���o4M�ޭ��Ow��9�M�ݲ��DW��#�Ύ֭k3�߰1�	��7-^��� ��M�� ����ċ;� � ��A�3!�23�߁}��\���Ո�ʄ���_�/�8��Y�8�� ��c<D���M�C0�3�~[�ua�%Ȥ�����Q��ȹwf:�e��4Sr�(׬m�c�=���:̟w1�$KrJ�����ӓF��j<��X�b5��9�?�l�U{�h�tG������,��YtttᲷ���z�I�O*�	�ְ���lX�>�c��/:��=�D�˅�D2�@$
�$�r�0��V<��X�v=��0	g�5��N��R�9b��~?��\���6�����~�aÚpڜ��:�� �RK��y�Ɲ��_1>�c6mڂ����8�sp��Lw�Ͼ/��K��{'��!�z,_�
�?��<�TL;a<ry���A��qə��4��wo
-z��.k=
��rZA�V��>�����Q�>�W�J%�����X)ۇ��~T�W�5�D��/Z[M�a;����wYV��X/�y�[�����N�3@W��5+���s��!d3�\��l ]�Y��E|埾�`�ʺ����?�굫LY�{�/�������@d���#F��|��e\��n��4�8 ����TPƢ����[�+D�qs��x
n��F����n/�2������6,\��x����9g��{�5��m�L+@���[�l���c�+8?�@)n�]���Z�3�8�=g6��X,�7��#�4ͬ�1�7RÆ�Y�ޓ£���T2��_~b�r�����ϥ�Q2߶T+^Y���|��:\�ˬ�]u. O͛�T
�]J��F��ú�m�5�$?}�{}�s'���'�s�JK>C|o����i\z�h���=�����/C6�|�e�h۰�-�*��r��"�NWe�u�.����g�o7���X��q�_�f.�c��|�k�1�KQ�b1��N��f:+5�?���w���0�1�r�-K�.'
�_v�"	 �>֮Y�|��~�N�Z��;����Rx�o�G�2�=�|�
K��h�������cǘ_��DP�G�>�y�|��?Sx���ٓ��E�ބ�e0��;�̨W����װ�����J�+�{*��
��J�KqM�'�?�f�2w�ҥK�eFk��t٩����i����	ذa�~�^�7�����/ K~.�zC�wc��G�c[5����'>���aX�n#~{�-�M���R��b�����A��e �`J�>������z��]x���8rT���]�{M������љ�捛�i��j/����5r�Pkb^��f�?>^y�#l���W��c�a��ٸ��������M �8L�
�-i�}��p���bx��U��3�.�ɓ�@0�u�UV.����o �?ņ�x�ѥ�z�;.B4l��������X�ڳӹ(~0E�P����.A(\�K.��/�p���L��.64<�ebVK��۫�x�_�~�F��'Ok���"M"/�P[_�\&��D���5�"�L��������s�%� VC-�Yg�nT�� ��a�0RE��*{��X���3;����ٵ˄K0A6�<�����ۑ�&QS]o.��x�<�֬^�Y��a��V���teutbյ��l7������*��;���=6�����OPW?��2�v�4����~��]���?`ƌ�s�$:��]�1���z�5$)+��T�a�O��4������ǌBw��(��6!���+�D��h�hG
�0v�N��+���E.�L(�]q_��G�sޥ��@�k�B��ʖ7[HnQ���������R;ŧ�=̿�׮]kץ��Һ�3�O}]�~�>�.��`ێ-�%M7�ջ�CX��{�ص���}�1���Z�v�e����^�=o��/5J3�|>\r�[p�y� �����e�b������2��>�5u���@ۖ����_�N���~��X掸��կb���fR�8����$��1����shp�H�e��.�/ҫ����`��-XH��gҤ1Ȧ]Jlk��6����G�Y��w�!W̠:V��;�X��Id3�u�y�U�H�hEZ��Z1z�K�?�^�;�	�PUU��k���Ï���W]�6�	�|Y�=b�}�Q�ݳq�F�m���mZT8T���[�5k�aΙ�b��#-x�L ��Mhmn�豣-��qs6nX_���~�b��O��@����CJ8A���    IDAT�������l��=;�m�f�X��b�Mx��'��P�K.���_,�b�w��13z��֯{�V�������I�m؄�'LŌ����k���c�����Ƙb�q����B(�@���������a�Y3��\gV�)�5c��񨮪Ǯ]۱e�Z���.�T�~�I1k��Y�`ֵ�y�9��˦����-��=Q��]V���Ą�c�򣻫Ú��6��@g�[�m�Ν��L'	נ=��,B<�,k�ƛS*D�AyU�W���ڂ��H����}����?|_i��!�s�e���[�j�^V��|��!�
N?�t�T�g:�n�Kصs��@���Hg3�ҫ�fV�K/�6���W����܉��.,\�PO�Y���P�oni��������1�A��uj����x�ϓ���ш�n� ���ȫ=��>�4^X��Ip"���>� N�}:&N>U�l����I+A�L�d03D���>6u��0b�H�[�� h@����ޟ\DFJ��~>ܜX�:m�����X��l���w�-s���I��M��L<u�����8ַ����]����)�w�"��_�֋�P��a��5b�䩨�kp�7�70f�<�ϊWV�i�}�jq��������Ǝ3�j��Tr�Y�ʺ��I�i�},��U�0��,;)[�"�ǔ��[u'��\N�֬Ya��-�:;�x聧lc�����\�8��駝�|�o�[ca�%��3O����m�_�����!�O�=Z�����Fw"oEl�\�����+m�؋a��Eذn=fΚ��'M7৛�����8�����b):�v#��Buu=~��[��쬳g�e�0d30�9u��o��@8��ӆ�<i�Z���W�5n���'L7Z�L>�qG���e�3Q�*ڸa-6o]i� �b/,{�=�8�;�\L�t����Ģ�8y*��u.���GWW�7;:��ol.|�l����c�1ۗ�1�_�ֳ��c�o��,)b^k��\KS�Y����T\��ϸ�<�v*�&����F��شq=�a	6mjC!�A�u�˙�Hkw���8��3�٦r�=��w��]�v�ǧ��?����"���l�5uHuw�8���p�EZ��ݝX��9�̙����S�Zpgډ3�3���n�����ؼys��YY���������"�b�Y��O�w���\D��SS؟�}��I*Me����ތ �s�������QG�1�3���N9���
w�옝ǚ�+L㣏���E�6��[�z	jc�( �#F�ńc�������*dy�]���=F����ex������dc˴A�-��`�6ړD%ScGb/���æI�U7�~���u�}�Id#�5���N2_��9f�6+W���V��Dx���gA̿�\��ģ"N:�TD���,hcЕDy��6�>��ۆ����g�Gĳi��@um���#�M�,_�ľ�Фe�K/c�ɳp�qS-B��ة���[���֬{ъ�BA����n�bU8�hh"wL#F�������+���M'���{v�et�btIΜ9�O8��+hI� qԨ#��A�H8�]�����9 ��^Y�Gys,�j2��4Z��q��i���?B.��/����L(�^��>�{v�j���z�`���_��_���Z�5n��3���֯ ��?�9ۧ�����I�?+������bP����n�E*k֬r�D��{��ZP��9s�c���1�-��H$q��oǣ�>�)�Km��A��@�@>��?v�����;�\ǟR*n!�15 ��ј-�Ԁ;w�4ʆ�^z��wS..��'L�����7e���5�QV
NБ/Q!�����ӹZ��)!3��4o��g��|s瞅Y3N,q��L�oji��ˏ��V%�k�V�?����Y�=�l=�HG��Bc�(TU�ώ���S(����c1m7�{���G�Ōf��u����BC�00W���8R(sh߻�,��K^�Ë�9���̓���n��I4Է���,1��Mw�5�hߍ��^k�I@۾5�+��#��3�c?u���kh1����WU��u[����2�}̽�|�9�]{m\he�@2�t�w�EZ��oCw�?��ο�0a�DTW� ��Y�OK�&�
E�2L�d�;en#V���;�c[.�w	F��6�U8X���ᨎ58�K��H,׍ή=�h��K/��SO=m�o޼y���2¶P���Z˰���u�T�,���N��)�w�h۸��c�%f�dShj�Z�2;���YDcUH&��s��3	�}���a�fd�yK�e�?W����wߌ#������Be�y}��3%RhP�E�u��FL�"�Db��(����V�y睇�有h�4�R�o7� �G���R>I���Ltw㩿>a�E,2WR�׸�J������7���OM"��t�3�	J�?�S�֙��,���0�E��1N	ݨ��}��f�o,�Rր5����rQ0����9MEf�9��/e��g���(��L�C�|&n
ˮ�pՕW����@w�����K>Q�.�?�����"���M��M7b��H���e�����;j�Q�2�̾����sK�����_8��0�����d-��M3E.gi�N�8Ͷ�{���m�މ�-Ɨ��O�h�oFu55_f� ��U�1��&�Gx��'��_�����U��,!�\��L��0��-%0_�r���
��w?��O8��Ӎ��2_��1�ч`�u�rM;�&���g?�)V�Y���w-&M9�h�K�D��'��j*(X��	��꘽c&�ړ#F� �l�s�C,,еBM<C-�� 
�<>���z�U��{fO�n�,��9��S���4r��ձ�(���o`��Mx���c��wOյ5�˰��DB��,��*�4���;��o�4Z#�DM(H�z��yy����ތ�5��M��%���ܫ���-���ζ�<���x.����*c��!Z�sΞ��g�RBp�%����?T���1�F��G{�^hB��6���"��ń[r�z�5���T�~��@.�\�}�J��Hu'��@��#�iy��H�B]��n�fA�%K��ɕo^t�ܨ��\X��9������^z)���
�F�lق���[#��G���V�'`k�_����T�.����@�wް����ry\~����>�qJ��aʣ�8�'�p���6[�KKK�}�{1bdS)>�F����N�s��r���x啗��}����y�7o�c�$�u5+����L�|2���p����w[�ͧ?��3
���8��
8*
Z�Jv�>�X˖?�[n��=i|�_G��<�d(�ppEZ�7[�TM����p�w��{�ԩ���>`<F2jst�T�/�\�b������ ���obÆux���o-6	�|_'����	���eEV�`���}�߬0�C� �Zb�V��#���F,G�P$%C�����L%3֓��ʀ廮yg	 E]"��3��T�Θ�
�mNw�܍y�.��g�m��9����UE1˭�.|�_0��B|?Ο���[kwO/�����@� �G�2)OR����`���c	�7\w=�=�XK���c���5��Y�O���B���U[[o�>y�dL�t&M�d������L�,e���|�)l޲�h������
sO��7���6s鳙��L�&��<S�"�*�U'�{���䗮.�<�6,w��=V���=��w��]��f�� �3������q�@�[�8�>��{�\^��3��mWX���9�b�JI�GkJ��|7f8�}p�u�YIw�l��Vk�n�Oƍ�ϲ����o��/�%��s�W}�@��>��������+�.�m��vwZ��EpV���Kˍ�+�̚�B���j�g̜%��	aG����\�Ɍ�p��Ԟ%�պ��b�����������1���q��e���]�������|�Q�Z]���C�z(�'Y���*3o�k��S�rt����OBC6N��Hi�^0�k�87]ݝ��׿n�T�gS�S��"�ý��<^~ �oޗA]���7�lV(Ӻ�}*��r�������q�l>}.�G����ɬu� ��i.g�K�?:W�cj���|�u�p����-U�
�mQ�g��"���MWcN�?��?`Ŋ��;0q�D|�S��2m�iS�I��r�G=L�mj.Ϋ�~��x���ֳ�y�6І��o|Ê\�r:z���p��ӜB�*�a��͂\��R߄J������c�Y����3�\ݻ�F��X����.!��\Ι�Ȕ�}�=����fw��ח����	Ǣ���^承���5�	��ZR%�/p�W��SL���8{�7���\s>yi��p��'�ۇ
�2U*���;�k��`3�>[~WIx����S���]��z���>��h^��Ũ�A��aP�B���O��O��3œn^
5�mR0+�G�}�kMy�0SkC�$כ�޵��$ �����n�����������p�X������<����޻��x9�,��O�Q:���X��O~?��O��SO�F�R���9ܸ�ٕ������fk���ݍ�����J�����GW"� �]�����C�5�����0p!�s�y��>�7�s��Z��2��k�E���6��s��eQ�gq75�)U��[g��q����,S榛n*[w^��2}J\�|>+7�O�Ss��M�Vp���y���l�|^*�&�k��XI��k��(tLP��Ҝ�7�T|f��_ti��#KV��+i��%�3��?�߁������@��>��WZ��?Z����g̭C�g̎���ts�QY���s��ˊ�Kq�
Y�"y�>�?�'&X��N�﷍�~�Cop�?4��c5��4�}ьg�We�X�/�R�����4N��J��1�!^��z\�W_��JD�'�A�K.
�?�;Ǉ���$p]{��S`���ečB<���E4�p"ë4 �ݧ)N���}�ƍ+��qC����H��y�	��ɭ�}n�� �����bޗ�?��,i���:+Ҳ��$���
��j�^W�B�"AR)�J๪ %�����r���T��S�j���eM�	{^�;��	׃,!��[�x��i��)P�Q��?;����˕ƹR�W
��k����ה�s|��x�	k�Ƚa�%>�]�F���ԓf�U~dux��!���h�aY =-��&m�m����F$['9��`�� B��w�X�e!�}��ɟo��?�ϟ`Lp��T�s��I2���N���DN�����G���l�C!z��� ;P7[������U_U�����X�?�~��_ۦ%��%����njC͟�d�,�� .2�ļ����PY�CAI��c���3��4Tj�^�qf��`�K�}��Oa���,��֟���1.fi=��~��aM�XZ���������{���l�e��ɱ&s's�Y��:��)��b�.!�w~�N�JH��Y��_�u�[��������i��X�g8���?�b�0��H>����%U/�MB��� �<=���^ӫ����ͮ�+�Y�\���,t��(��뀚i���$�q�8�Y%*��1��]�a,���{��/~Ѵ4�T��Wr2�-G��[���	qik�*cD�A�=5�z�i�H
��n.��el��.����O�����e9h2t7�閠��?��Σ�e@� F0�Ї>�Oo�Jc��p'��y�FL%Gn����z!�݀�g�u�i<^�Z=�i�󹔦���5ſq�8�|g�>�@�8	2�Ko7��u貚z ^kDs�U<��z���޷T�{��������������$ؗ�X���:�O_2����4.
Uj�	�<N��?hr�?�k�߻�}B��]���]�8��N	�D�f�]�L��ޚ?��c�l+1��tKP�_J�/95p�ɾ�8���ÏW���ڠ��㩽3�[�L#R����I��k��V��S�3�ր����o��4L��ILŀ<0������7O<����]և��g���g�	c+�w�
����TO�+��FA�Ɨ�Qh0���)Gj�{��eE����_��=��y����j�e���d�p�6�;� �  -J�,еT]O���'MS8#�����/,p-y*���#����;��������.kS��ڽ7��w��˔���X  AN��Û�9�f��	��
�)�h��)��{z�!����� <� ����W�}�9�=�I�A	������[np
 �'��&�O�;��;��\��'�+��c$���}	� ��Z��b�6Xa�M���!��@�^�KS�'S>ǅk�V����/�嫴Β�q �+~�ؐ��v����x+��9�Z���)�%O�'!�w�6�h�Z���s ����pK�'ô!�D���+�Sօ6�ib%��-��e�-�|���8-N<���� @@��`/^ %ׁ�&z�M8������;�_�`����C'�D��Sȹ�G����0G�����	D�M
�@�a�����5���xǍ�4i�;�8N�|x�� �%Ùw����j��O�^vdJ�q������'��&L���H�Ф�4���Y�}h�|@#0�4\�+�b�=M|P:�,EU��v�.���T��J�r���6��L-���W�Cg�qo�NU�e�Τ'P3pK�?�2Y��L��1����5}Q�������a�)x�
�x�J��\�C=4C#``�(�}/�v� ���<NBA^�O��z]���zPk��R:����'Y�7ρ�Ţ8�9V� �	�B�-غu;�[�Ě�����M�''�Z�R�zg�ȊP�N�ƿs�9���|��ch��#P)���׊�oJɕ�/OS��3L`�8@a�:��޲�z\�.�Hx1�����r�m����W�]��C{�O7P'�t��'������3&FNYɛ�((Ĭ���>���◿�\r~Om��}s)E�o� �<�N�1���+��Ga�
C#04o�(LռJ�^��8a�8��!y��*Ͻi���1]�B����Ć�ͨ��`/��^{<��J>�P�eeĢ�_��y��s�8[�������	bfN9���햮&>
o~/'�����=�R\4��L�!�#���=�F�Ў �CY@��`vi0�2�|������V�R^�J�
짟~��՛��lP������nG{�#���2诧����_lz-M��7m�|���Y:#'���	��g�2.wJ_�U2��Yy*�~
^�a<��y�����GB7Ѿz��eedV�e:t��������U+ �Y���8�����U�KE��_��f:,DzH'���Xu-�i�4�J#0o���������3�k��Ϩ>����4�]��h����O?�-�6��C���c��)�����z���D�NV�R2쯺�*+���?h�b� ����}R<f�7o�;5~��Z\�P����8�#0P���7
�*������pԘ��
ho߃��_���/�9�$4�c��4u
N�>�N�2X���F&�c��{v��;��U�b����>_|!�?���GG�.lټ+W,C���+״�]��/��a��=hj��_��r�.��S*��6"�<�<I�JA@:���;����Yu$�>��
)�W��C�d���f�J��ߦ����o����ys�	�T��=���d��*b|�ᇍ+I-���,���=�C�,V���z\'������L��p(�DW�v�1i�4�{�\�&�F���� 	#��b��f'����y�e�+��6K�[�p��cxk3�a/�#G�!ѵ;wnF"�i���c��{W'��rؾ'���0>Jb6V�_�B�yK���ok���3 i�#�7}�C�."c%3�xi�io�3�t:C��#vx�W���2�L��� ���q�����yZ���v�a�
;�>NN+z��n�_���N��X�a!��g�KN6�ö�q$ytv�p���4������� V?��R:iI^�7�������s�W�y    IDATq��{�����
�|�tn���s�I�6)������=�شq;
�0�m�c�)s���Et���R N�.R�ra0����[p�h��j����xQD��t�!���n�7�Շ���5+^��N�\�l\3��#ͺ��ץ�;*rO�Y�7��Q9���?���[:gW�<���3��uQ�X�"
�����](ॗס��	�mÉ�N�o�d�ܼu�%�l۲���{�J.�\sK�����m��o������!��z�أ�~���nj[���g�9�|7�n_�L*iڸ?@n�6�����6�cܸ�֞Q��_���)[L�z�[�b@O���"sz��E�����:(�;yq���(��\��o�i����5��`P6�ܲT����O>e��dOe"��(���iՋ?�$}TIHw�S�ߋ���ں6mZ��nrd�ΐD2��ϯB0P�ݻ��|���~�2|�E?��f�Y���D^E���������f{{���}�l�Q��cƖ��W��p�ٳ�Iw`���Hg%��:;��~�&�|�X�������C�`o�(jt��[]T�Ϲe���i���L���RJ�����������P(�����P=�`��hY�1N\<ܣl���6�ai��ʑ���I��fNl]��Mvu�����˟��܃N����jlܸ�{��J��o+WmD6�Ggg;v����/C�%�o��k�������#�Jc��1����4��R�N�~��p֜���Ѷq5�.͓����q�m؂L&�u�:p�)g�{��y���;��'�D3��6w����L�`�L��9*4Sw�����{���{��4������¡r���_��/��]~�=Nk�,����~���]�� ��><f��x|�]�4i4ZZ�a��W�˧��`c�4��+���Ua���5���n�����;�������imn���n�y����������-�i>��`dK3��<^� F�jB�Ѝ�{�!���y}~?��3ؾmv�N`��$\�vK�$�3��\4�.�"q���ӭC�9�	�����;	�n��~�LM>���c��^�(��}�ڱQ��.��7~�������;�q�W�ޥb���g�q����E�̚�`i�3`���]X��"�TPc�捌��G���;;�ص�\x	�=�D�bx��p�-�X:���+e�Z��/ۇk��<A6
a޼K,�3�Ma�m��ٻ{��B��k��<�gG�6lC8ڈ��q�;'��o�TOQ=|�k_3�gF�z2ݓ�AGaB���~`1 /{���6���A�zd�܇�y�ߐ� ,�_���"�̦3�\bꕀPU.��ty��M7�d�B�5l۲{vmEGG;�9�����l�p��֬݀t*�+���ǌ����nK!��������o�����?P�o��#�3a�x��w!	��&���������Ĉ������Z1�ē���	��g������ގ���:�������N�nQ{V������K�ސU���uoٹ����j@��U�C�痦"�h/Į��^'KJǊ�[)�bB��\����MT0���(�v��y������y}��N[��Z�I[Ԇ��[���?�2AҎ�W�H(��TO+D�5��i�0F���K�E(��3a
O�/�@L����;��{Cc�&6�{;�ʚ�R�����uEE�)�j�#�@֬�-���zy8��_����g�{S{ϻ�1��w�m��T\T��I��S3"V�~���<��/�͛6��/����ծ�u*�A8�$S̘q2�u����mہ��zK3�{�R����y��?���R�7��ۀs���ݍk��N\tх��E0�����F�����{�PX���b�'a��3W����R5YuG��6	]=��ԧ,��_�2��f�i�`ж��|Ŭ��������ڜ��`�^���q1�	U`L�`p�L��t}��4����м.c*e8H#���ܔ]t\3���@J B�,��+}O�ϟJ���Ϟ=��*�CA}�(K���^>�hx{[r��#�c����	�us��GY�p��[Q>��_i���t�h<ԉ�?���ΝkkQ���i}�ƍ��̵*^)i�<O���֐�U�\o-���i��IF6Ї�s�g��SO-�K՜j\U��yb�<��wT��~��`��E�G�/�������'5s�?���bʔ)`;L�'A�}�9�=ʣ�c�����D�f�j���{�j�
[�&p�>���KQ_7d#(|����Z��b��c�����h�hR6g)V�lʢ�'N�n�܈�H��,��0�� ��"",��Հs۶mX�x�i��(h+ �����җ�d������Y���H���j=��{��*Ս ��w�۞�@��'P��gg��-p<�
��g�8Â�
��$�%W��o��o6�2��o�G$�]w�mD�e��w�	�����a��s$�x�)���i�eG3��T�Y)ܴ|Ư��e롯���~̸��n�^��nu�i~>�����M���c�# w�R$�2��*�'����-�%�sK�X�I�����2��J�*�4Shm{�y9�V����&��@��~�T 4�R~x-u�b^�O<a>u�[i��`�`�x��kM��t�R�df�=�̳x��l���
�����[��_��_mdAr<�'��'L��"�t⬝R��'.f���/��K+�;�S(�����/�ws<�q}%�_Ҝ�C!ׄ��/���/�	<j�X+��ĤS�=��ng�Z�Ҹz�z�ro�>���M���}C��Y=�<�pT��i��]o��4�ú���4<��;��P�������*�Z
L��XȦM���8�K����c��/8.�P�|�[߲":�6��κ�����y��n���sx��|�,
�����YL,ܡ�ƹ�Vʟ�'���P�'����:Ӧ5!W�c�����'>�ѣ� ݝt�鴍g>Wj���~�,zx12� ��"��&���4�\c}��$׮_��~�����3�
	�a�?�S����Ϳ��q�1��nPo�y_뀱�5ZT�����߼�M�b�}T����*;�DkF��K�Fp_�z��w�'�t*z,� `��:�ݏϨ����;�-�<y2����@��2�@��d&��h���x�������y���*��d�m�w���?�wį���<�M��/���b	���aĈQ&�#W��c�m�b�H\\�r���2k�,�`����	&4��{���{����a ���X��k��|j!��%���9K}-��	[�)]e%u��i����oV��y�j�/^���{���J_ڧ�Ҕ)|9����%
�4�e�!����q�Hx	�5��X 3�.����b4�K^��||^��8j��}w/��9�т��z;Ə��ꪘi�Ŝ�1A�߬�l��N��~�%K���b96����80퐂����y]�?߉���_X�̲�<<_��֯\�\���ϟ���>�ƕ��j>��y���J»�:��B�2d8��I(��k�YY@�5 k�d�RYܡ��^UV�u׾����rl���%v����*� ���SӦ��jL�:3N�i����Z�\�(�
ؽ{�Y�_|˖/�`�Yxp��IH�ߧX,f�[Zo���^6�����W�` l����h;%-?2���}���b�č� 087�|y\�
Ԋ�� C�+]�r��Փ��:s�L+�b�@n-�}�C=4K���"?�Lpj`|~� ��ǟ\���h�`z%�g������ K��UV�5k
��AG�$�;��I��97��xg�mJ����^ם�W�����1�t������T\O�J��}!�PЇ�G�D,Ze׬��3��s���Z�w2�l=���� 	���"1#���lr����u(5>r7�
'6$Rq��Fg/�*�D����1�y�ǖ ���WZyA��N��8����\^|^^��*/[��x���Z��ť�����.Ɯ9s��X������~r�0�DE���U# ˓���pMM-fgry
��)���q�;�]��/ 
�?�p�T_�Kk�����{��_d�h���v6n�w��:l��6`�~̂�a�	|4u��5�F޹���h\,��c0�~UnP��e��dpL����IVgi[�78d�3���M��Lݔ����H3���+�?e-�R��@����~�^KMA`>���	�y�,+l���u��y׊e����r!�{�����5�.���u�}|��<�"Zʱs�Nz|���[��Cw:�T&mY�W�;m��#����!!dq-�)�l�("UQ*~'A�FD;�#���Z�^7��-ŀ�:Ї�?݈��y��'��\^��)6����-�,^�1�Ә�8a�Cʅ�C9�P�"�����82�ɖ�,�8]|ʝ����&L�0wkIY�4�C�_I�/2G��l	���}6�����28_A �w� ~�}9�o�<��XNjE�C�'5f|����P������O��@��p}/_����ƔF#w��@��m�k�C��8�jb�ո�	�x/�W���'���=�Q�,�L��|yms[T����+뽏6�4P��xm���_
Z(���x�Q�o?y}9㓊R������w3Ѐ�(|�XЕL"�ݍ��%BB>�57|F>��G�{��=��Wf�U��?�nP�}Ya��������;�0J���T�Lk��O�TP_{�{}	cY\����|?zo)�^+���|q�r��w���|���:�ڰ���,Θ���w�Wpk���ܰ�C�8>-�XUM)�9�B�Y���ks�u����@n��>���Uޏ_q%߾>��O����j>.�o~�.�\^��b�t�wmmm��HM�	�|z�q�ۥ�b����w>������c�F���8&qӊ�n|����&PB�2���9����
��	��1�j�����	_�ц�������]6P_�� �E#`?	�;ݎ��,A�� ��է2�}��V�[��|pL-1@<��2�4~���ZEWy�5�׼{�Mq�}
��ރ�Y�W�e-����y���t��Zpoփ�8�R�O��SƞR_��y�A���[0�g�xǵ�|�}�������k�k���11��c��w �G�r��R��w����'�&��f���iԇ�k���m����*ȕ4z�p��#����������Q;��W�ل�G �{�B	�$ zP��i7�_6�����{+��9���WC�����aN��{�B���L!fŰBPy��'�Ng|mK�������b�U��S�0���@�����;�C��k����iT����*��c=އ!Ϳ�ٚ�`�/�����^�/W�4x�b�?X
ZQ�C�!�]�J���K�0y}d�݆����}�f=�s�ұ\��E2�EE��"X6Iݜ���S^�}	�y]� �==ǻ�D>�5��o<�~Me��_�����p�L���h{�Y���8��K�;�w�Cm^��R�@~�ײ��!�?����>N���t���b)�3�C� ���>�`	&�B5����|�S!69���A�?�~_�P�˗�*X�0�$ �R�	�S�2�5��e_4����!�?|��/*��}z�?��l���3�K�O#������p.������e�x����W
��J@����A��3o@Ϳ�p9��.�n�G� C����uL_i}"�� P���ؕ�/����^�UX�C����:ʜ�ޚ����3��f���r�i�o�n9�{[O<z>����{�!�<���_(��1��7����qzh�;I�$	 �M)�._7d.Vs*7��+����a��}\@]�CK����+�?}��Z:�?h�>ݩ��;P�t�!�?p�}�a½�z����U1�� ��-����[���om��`��-X���x��*���A��9_�:���W1o��0&�������h
�L.�M��������G#~�@��+Ư"Q7�U���U,���7j(e�0E���������"P�~��������ZB���R�?��q�|t�Z<��*�Qі\i,2�Y6W��Ze����y.�->�ݔ���1�G�����0�^�z-C�S E�9s�(�O�U9����nx�p�d7�錍m&�~P	QV�����|V�6���J�9Q"��p��*k��s<ʬ��b�bU^
�ǎ���X�� �k<�TZSz{+�5��ޞ���Y�益=�{C�Z�'�jo�^Q���G�\�-aV\>_N�渲��\=~ �h����=v�+N̻b�e˞7�qWp6��?��y�"���������q�?W��E.m?F�����zm���>V�=�B!���&-�j`�&K��k�8��*�i���#��?��% T0t8��\�L	�ci���w������n,��R+T��Whv�L�6���U9����K'皙x+O�!is�oW8�tm`iS(�"/���=^��J�������E�+$^���������r�����@��)巪^�hir�Q�H��.9��8q���lh̩�X�TI��
�%�����sz]���~����|g��8�t�QPp���sq�xoS�I��kk]��������)o�s/�'��Ϥ�=�i�ڐ��U��.\GV�۝Fsc�1�2|ذ$Sd�u䆉�k��V�$�[���9\�\M<�p���/��m,G�Jt9���g�y.�{>��r�O:�4nFiuiv_�۷�4C
m i*� "��F!�	���w/�x�B�`��F"�i�RW�~��/�1I�Tۻ��	��	V��x��}P���N�J�7 ���#F�w��W��ss.�R)mb�8���;����x
x�Yc-�d667�S��ל���_ȣ:Ve�.���pu �Q4��
"�c���Y.���������:3-��E�,&	6�#��(���	N	X�{�ݏs�{h�Er�k�;����Ha�߇�E��,-	j��Ƿ��ގ�=^
/��'��s%���g���0�Z���ӊ>aډ�����W�.�h4�ؾ�:s���T�zV�X���q�Q��-�@�ɞ���/����x��>�>$v�3kcU��e�I3��oKS#2���X��Yk�F�-.��ԩS1i���k���.l�B�a.|.n�#�<�ƍ3ӍVB���M$-�C�?�:��~ ��MWGg���h��_<�V�	ۻ����{r3�1������ �U�oV��m�L1	g��ZB��TE@o�W�KSK�Ϳ�CZ��xe�\�Qy���w|G�]���Z���ޝ�_Ȥ��҄=#���]���=w����!��RG����f-!���Xr\ml
���:+a*ˇ���J�)	yZd^b;���8n|w�I�=	��LyǕ�	]�	bY�K�P�{o�Y�)���:֫��~N�:�����~�s����r��9%(�F���q�U{đ�DB�fRض};�y�i�w��Z�Ţ��;|�H{�h�Ŀ�?��'k�h�i n�A����a<�qc�oմ����q��ދ�G����(���c�`˖Mf��������Gy��v2b���nH�L�~�7qQ���<�_c�@n"i�2����5�v�����˟1o�E��H���|�I<��2[%��ߩu^xᅶ���
8R+	@���&�Q�)���x��)�i���8q�]OZ�W�P�}�=�II���^b.�#�l�C�^j���e��r�xP�����;y�P��B-͍��c�8��+7倾�]1�<y�]w݅�/�����F&H��ƙk��#8_����[��yK_x�>�h��D+�q�e��36GlIK^S�7ޗ�p�w�y�)Di�_��O9���J4^��uE�C6���l�Ə,$�}8FrG��ټEc��,Y�[n��L�,�X<F���1a�8�
i��	,~)^Y���&0�!\g��L���3g[G&<��_����j��F^\�7�s���?h��?�'�S�.����w酸���+f�N%�f��xa��,(GL�O-lW{J��s    IDAT��������r�����F�L'����6�}�Y�[��� �!7�c�=f���J�����;�k{�K�5Ea�9�6��K�$���{���\m�����5�\c��X�x�cC3�{��6m�\�*�F�v+-��8y�d�i�r+�Y�.
�qd�1���K�N�/�7�bw,cW,���s����c�<�쬪��N���IH!	%4�]P��2"��"
D�*���S��\D)6H �t, ��i�L&m2s��~������̙3%���'�̜����~������Q���ި a��}6��{�=���FΪ�j�p�~����4Z>��#�;�����f���Bs�8���2^��/Y�T[.ug��Y�|G�\g�64���˵��|3~uS��ڧ��ֲ�Ro��#���4S�Y����9R��q{)��T�E<�|����i�(Bt�y;J��J>�!y�'���u��qo(�\p��Cy�S��?����V��{
��"�3�.���mr��G��%y��X��t��Z	8���e$��� �l�Pe�w�o&��^q��2k��2]��c�� i@���Δ��6Y�r��tw���<��w&,�ΐ�9�<6��p�X�[@�Əf��~�i�%Lb����!|m�r�є�i�����y�W�blsr���qPbl�{u_ɺ1��5`��f7���D�E	��ۢ+��h�ԼV��i��9�����g��5��� �W~�����C�h۠F{�6|(���i9h� �O`�`lX�?��������t���K/��ӧ�����k�W� *��oֱ�/���	L���s�Ygi�l���1�e�*T��9��́�N�lNۏ�X9�kZ��0��DkHU���|�u�i���|��k�T�� �Fu۫~�k�g�ش{�=���|E׽�]�y��=~?��hw{>�=~�}③ll^,�T�������˜#�X�(/��5M�$���u媫>&3g�.�lA�x�or�=�H,��}n};#]��~[2��J�j�O�� ���ڨ�}�r�����r�rI��f-�M�NGd��9��cK}h�������	�S����Р��CM��S���3��r�����8E��̵r���1c�>����#o�q��hO �i{h~F�������K��u�P7���q�  |��6W�k��J1�b�?�^54f�Q������yJ4E��q��&(��Z�v���_j�E����瞳w�/�P��t����E8��Tł������ G�q^�*��;�MPs ���35�ߴ}s�+�Qp�6��)SJ��	_w�y�j��h��Dw���t6�6׀?=|�^0��7ø�m��+��_���9��W���UysچR���i���ӟ�eie�yN�w��Hn�g�zHƍ�˸	�d����U��tN�-]-�\X:�S�����sϒQc��ˋ^����_��͙;��ɶ�+�?�3,�ٻ�&W_�!���ic�<���r�GK>�%MkWIgW�ĢԨ��斤4�k�l6&���d���Ҳ����җ���'�E�hٴ,$۴��'NP�0-�4EӺ�Kܞ��s����cƨ�vb �wM�t�E��pԨ�ȖIH�ײV���h�f�"�\ )���`416\_Z�?�/�B�'�d=�����E��s~��|l�an�]��/��8-LШjh �1�t���CF��o�k��8�]��q2f�o�ͥY<G��9}���ic�o��8KN�~�X���J�w��-��x�W��u{��W��c���uO�ߡ�� ;��{��gk羦&GU�u��O|B��|�+�'#���3F�,}��ڰ'��c����"�iiMI,Q/����$D�I.�ma0{��l���G��?g��&����G��s���#WX"�����By�O�!��-�XA֬]�m1�
��l��.�6�O�F^^�V=�(�B�(,P8bQ$��pL�����Xx�Y4A5����4__s5A��-n�O7��1�	Rv^�����67	b�e���>��kn}�ôG]��xWz�:��1���� b�c�����>����S>���'��ρ%,q�\�:��U>��/�?��aB����� >���O�z�{3Kz{��Ӭu��>�\N#�h�������{�.8}�~��l}A�]q�J�-_��<��{�G�'Ə����)Ţ�ĥ�+/˗5)�l��)�Z;��o�Pԅ��䎟Ȋe�J}�s[�����j�Oz5u�NS��k>.�b^��.��m��c�L�]6nZ+�=�.����d�4��$�y�ؒ��{�E���*~4>�i4`�J�^8M8P�p���;��1���Ȩ��6y{.�j�f��Z�@�`*�8L�y��}��7�EE��iަ���>3���=�����;����Aɿ�	=�,�����ܒ���(�&����k�v.��]���+ 6���o�3��M �
�	�Jc���߿��*�����s�������2����� ������Ϗh(�2���X�PfX(��׭�'{P޲�,i�8ZV�y]2� ?#��lFd�+�K$Z/�YIeC��]'��Uo��fY�b����R�Ap�������i��}��1r��?*�u52nL�,��Sy�>�J����u���ۥ�G�	i� �[��+#k�&��S標�Åޙ?~ɁH��SN9E��Ǎ�R��[nѰP��\t�F[����j��&f,o4�������L0��i���f��`?_�5'���K�F<�}4��9���h����(�Uic��H����l�|6�v�6�c�='��} �4�V�Uc��߿����)��l��������}'�/��y�fY�M���j�f�� ����9��w,,z_��X|��ΎM��ӏ�N�GI"�ի_�Tڕ�A{OO^^|a�D�d���r�ۏ�y��֤?��w/���������3�gvĂ�i�7~��-yU%ڇ�Y��Qrּyr�[����VI&7�����"�0 �➡~��Y׼Q�6o�T:$W|�*}`<�[o�U����׿��=1�h�\r���%�m���.�C��k	_��,zc�x8�/�\��4/_����/[���[>0�Z5�� ��7 �/��|喏��]������<>�җUe��K8�}k������J��ӷ<�}_Y�����6��/��p�z��Z�׵G~��7_�~"��?�|����͊�Ә��@���j����ѾQ2�N��R��C�����BL򹰼��5iK���^";�<SCA~�a���%��T��w��u�=w�}{����/���xC�=ye%�ϓ��T�n��v�X$������MR�Nm���K!�x�N�;�p�m�=�D7�勉ǂ��K������w����%���A9j��x㍚d�S_���y0���Q9�].��V3�r-��r@,�0 ���%`/&tʩ!Ӽ����W�����������2��}��\�3��e�F9��[ff��c����W����TK4�ݗou���r_�9�4}�����$`����Ja��l��K�'���p?����K.��2I��*���חȚ����t9k�#TN$��ttfd�Y��A���@$:.��^eFՎ���77�a�e��Ͽmā�$/�_#k�9�t֙g�	�'�I��Eem�Jy��G�E�4��E���C<DN8�d�0q���&����s>��'1���Q��	���-Ġ_w�u�v]�j˖-�gc��e��+4��6������26g_Ԑi���� �\s���G����1����s�F]�w}�5|����[�3��)��@����?._A(�r��`�mǚ 1N��90������1�[}��h?b�W ����XC�w�;\ߊ��Ӭs�s���WK�K�dlD�� ��<���}�{�+�|��c��j��_�����4�]��� ��g��M�9��s�}$�/j��G{T��կt�`�/pM����M��p����dā�����f���*���k�/��޲�d�i�0�����.kׯ�H$�^���Q�'���x�F�v{�-�76 ��,��,:�a4��{�q�>,6?m~��w�߷LO�2��6�m�j������V�7ЄmL�¡ڵ�|>�����7�-_p�S��P�Y۹lN�D2~8����1�9-⬿5�h�Z���i���ߟ�r���{���)�}�A���5���kв����w��cʬL���a��E5���:���.3w�x$*�|J�I(]�\-�J��<C����Db���勲x�k��L:���Ek)���;�~������)h	�?$17gyW���c�	z�n3R,��ڶ�X��H\6lؤ�(�`8{��q�<c
�>?1�"�.]*].�Ӿc��@o8����w�\����\��U��>ܱ�����w���	Z��\)�u[i>�\>������KHM8p.~�4q��}�9��{Hm]��pF�Ơ�s���W���ߟ����w�a�}/����
`���T؍	r�TzB�ϸ����d�ӴD ��<$.��W˚5k4-�� �Gc8�st!|�ߔw��r�W��C�_��7!�?����0��l���\~��-^~�9c��(�.�n�3���1��3P�ӱX |ƌ�g�$.�x�����߯`mt��[��:;z�V>��#d֮��J��m<�%�)����/��ؼ~�
����:�{�
��Xο��kRa�]c�b�uM@��3g�t��ٔ
2��E ��n�KI7��'�"c��D�|�T���p��iZ������V��b|4���YMPq�JiB���m5���1�n3`����ӸSj�S����Z�T�%�+�}OUU�^@�6|��h9�F���)Sd�3�&Ӓdv�x}�J� l�����ߜ���\�ol�)ٞ��R��{(��n�� ЇM���+�f�?U+�j�HfK�e�=��h��=���t ,�`���{�Z��~D~��ȢE�Jac`���l�d5�,�6����T���lc�{ ��ߎ�7��~f�PoW"���ֱ�O=�TU��A�ɜ��`��?�h��|�8w-��)���}��8��	ܾS�x9��jUϑ��6sa.�9����s�Ľ{ci�����a��s�2~��7��Q>�yv�Z�.b�����'�"ف<d���z�qu���ʬs��E�7i\���6�q��ގ�w�j��MX0C���Z�r������O�'�?��u3�9W�y�1\3 ^vL$���G��� ���w�+�F��?w���d���4<��SIO�>�$�o�]X[X ��kSP���9UM�дa���Z�2�V��pJ>x�AB"Na�},���!}����i�&��~�-.,�-��������������3��g_X2�%l�!��\����J)=y���{���U�H6�@�I8fmb�*KmM�*\q�Ǚ�^��M;�#B��#����xK�=yI%��|>� O{�z�Eh◭T��{�("�|o-u����� ��_ViM���a�QŐ���'�/�o�m�X��p��%�X}|?���E2X�J���p���;f��},`¢x�ꯖ=nܻM��('����5�q���Vp>�f:�v�D��������Wp/��\��B���,��3�4�������8�*�O�n,��F D� ~H�0���F�
���j�Y�u�c��'�.�����c�@����]�\��Ec��p7����#�4ݓ�s�Q?�EE(p,��M��Ꭳ��{�՜&D���1#��}y�m��a�zO)ʡ �bX����tc�z<7֓����	u��w���T�����g�r%,"N�{�iڼ i��^�Z�
7
��7�Is��G��d�?tE���\�4��
��.�;�R��Pi&�����c
"L�N2 ⺨9M\�GhX�
 ^V����
)dz%�����m�2�/+�ZB�{�k����Z�6���4�+>t����Pi)���L^���9��SUU_4�5Kry�21*E���D����x4��H��Hb���9��3���MH�<�Ũz���ϲ��֞�H��	�hB�Ǣa����ϥ�~�K졭g��o�˜�VEV�� yʀ�֥�_�)��o���xn�G�>2���
Ղ2S�d�}��P>4��!3�%�0.	���}O�\�v��sP�G6�W��#!��b��$1�,�6��� �Y�]X�E��D
���F�����-��s���?f�I'�K�w�y������ӱ�5	m��|J��X �>������n2�`&��8Z2y���$�1	�3�tHM�[:�֋d���HݨIR��%��c"9"������ϰ�Q	SS�%ߛ���l�N
Q�LT�y�Q+�ܲ^6nZ��^5-�C���~��d�`��VdN�.�ϱ+�3�����7!�X,��>��-�ʔ9W&ȸ�j���;����p��l�Y��`���9����0]��J�*�|���?�aҥ#��Ϗڒ��*i�L:@��C����a�e2���������g6�.Y�����r��6�Z�v�g�;K�O+8�
y��@�i��o���f��_��u����/
�c)�$ �m� u6��SN9I�<{���Qb##�IL2�uHw�
y��dݚ5���mǾSƌ�(�bA�E<�0�XC �<�
��Diբt��k$'��8I�k$��H1&ɶ6y�OԒ݉�:�Td���/p��̙��YT�$�Ȣ�,�k����O�����DùJ��	'����{�Z.e�s�b��}�����e>=��h��M(���zA�%��{4H�T+.PB��2A����_-��'~�i���k�FMM�F�(؇c[4Y/E�� �B�F���˼���n���P�M�I�Nш��e`<�̢��;��=)��Iy��h�#l��\;�l��Xb���!���*�l��J�G
R�I$�*��:���Ț�Kd����ݍg�����y���6�m��d�*Z�)���J6:^�?C�z���i�I�������vB��'�r�c�� @ȳ:�3�$	�>t�	&@��}[so���$f�(�ǀ�$
�q��aaS�B��������؀0N^��P= /�5��C�R?fQ���2�SJ�?��[]�o�4��YҹZUOʹ�)�ȡ���ۅ[9n������b��L������+�V�i�,Q*%�˨��F]�Z ��S)�ɤU��L�H���t���-5��&"�#t(
Ю	����{�±Z܊��D� �\���I"�"�^p�lްF� O>�Q����G�F���ry=����c�}$"�P��#�$/����-H}�hy�EjE�ui�x�s��{�� {Y�y��2�47'�>3���g�f ��Y�Ͼ�i�n��O"��XY��7�կ�ϱ��@ྍRV��r�Vp�ņr��ou����J#	8��ܵ���c����;��dۇ*�>,>�4��:�ҮA3�#�6���w�}4������
h"h&hZ<L4��1���M|���|�v��U���%�؈�	G$_�jr�Y/�x��82���wu���qN`C�`��c�f=|�J���*d�.���P��:W�}w�"��keڔ�2g��R;a���Tt�`�/�׹�)�~V�DX#��IE�J66Vr����b�F��H��I:�s�x�|U��P�7��8�h�Dv�\Y�4�ӟ������cL�5���&�:�,�����k������?�W�u8���-�����d���RS�ڻ����h�
���~�D\B&�SkE��׈�j�����N4�|XT�pL::�d��3��w��͘Q���1Rp��ާ�|w�,>�i4�%����Oߏ@���Q*��%w�_�K,'s&eD�D��gs8<��Y%C;@�0�H���p����3��)��&��i�f;%�k�����n���52i�$y׻eB�N��I�)��I<�W�@�O\�֑��|1,�P\ґ1��-    IDAT����Lx�d���
jRc��7|O��Z�B��r,�2��G{Qd2
 &<�֦�����G}���e�����G�{${�,n��u�ܹ��'��)K�B�ׯ�iJ�P�����Q=%� ��!��|��r�1����SU1����ē�* ��]J��T{�#��5p'�V�,׏�M���#o{�12��4M��f{4�C��_A('��P(��1��'�����vg��o�|���a����z��|Njh�I�i��pF�|�'`�!�i$'E�hS�lЧ ��n����@ ����,�^�7~�g��F!-�BJŤHO��������2m�t9餹�0e�tt[xja����POH�BB��h�9�	�M�j$����z�>C�߰a��薛�E/�0@�V�۞ c9! �瞫�}ӊx�-&h�ϛ��|� (�ƽX3h
�)��Q�*f{=#��L�(:m��ɹ眧U=�����&�F՗rn ����0�A::����ğ�T����j�/��dD�>��������G+�>x���h������|@b���]'==���+�i�Ji�h�D̳=��Kf�ds$m�f�7�t�.V���o}?���4����[5I�c~=�<��-�J��R���-?Q�?����Ȼ�}ݜ ~�����$���4�����w{�?��X]7��#��vi�u-ᨙ.��%^h�pz�ܿ��Ҳ�I�N�*'�|�����d�]D$L@��7�gP?�����? �/D%��tt�d��[/�P�&|��ٞ��������R�\���@��̔+��s���a�DЖO9�Ufx�[���<s�G��5i�ja�>�VC������k�[	��4t:pN�x��ަ�N3���e���I��J(pN�)@�˚�����YH�ͭ��ZP���=r,����#{��C-r�N�;Zeٲ%���0y��m�=eԘ��Jgg(�L��ؔG�Z.�F4��il�v�=��J����l&/ӧN���u���mw3v��\�T^~�yy�����E�A�%@gƴ�e�}���;Z(���z��'���]�t��g��P<���L^� <m��kl����a��5�7Ż��U	�K����$�RISP�����XM��p��%W�v���I1�)5�#��&��*���Ҳa�����O��:�cͻ0ϡ�4r)� ��>�� Ӝ�I&2�9|#��KǶX,!=]���?��!I�9�a8�>>�E��U�X8"d�J$�O���0��#�=��$�
eb˾cc亥���w;�ʐ�&K�4(,�p�PO4� }�#?��?��pn���_�Ĭ{�@Y�2������n�:�h��y���?��J;�C5�1�M��e��瞑�uM�A��tugd�]f�G-�춇��.��GV�m���9��w�?����B#jf��lZ
��,ym���ҳR(f�.�~�$�HWGJ:;3�����G��
��w��]u�(؄���g��?��j.<0u�i������g�yF��玚��x���P���L$H�l������m������s��(��P�S��Pf���[�e�j����j�)�?�揀��Z�B��֬Dk�P�JN�%������	��p�v�wȝ?��<�ğ�TW����۠% ����I�����wb�)*� D��c�t_����+Y`
ʶ�~�������������}�$Q��c��|���dJA�B�/0�J1�W'k&S����䢋��C�=�~g�)�����ַt�~tc����_�4l�����^��^]$�m%�^'��:I�����#�~�z��݋P��]?W_ k����0i�#2�s��9�J&�?^I�g�y_{����.�fH,"����"�F'��e��l^/==��$��rE�ܒ��%3r��)S�(x[M��i
\�f�Gu�nD��X��K��అl�}�-��K�`J����$�$ �A�
��)���}
P��JZl/��UMG���4v��%����������e'h�������0��|�o!\�"Ų$_�s�ђz�6qٸ~��z�O��?�4�m��e c`n`=����k����g�r�Ъ�<+V�(Պ1+´c�?h�"4��-4gֿi�f���l��QF	��Ϛ5���D׻��V>�����Y�k�>X����(c�D0�P�$��{�{�k_�����8���.�HA���p��4��/�X9�I�tHrs���6˺uM
�(A�C�>���^�^:���K�a�Nz����k�#�}�'ߑ�z���%���l~^�N����5��6�{���v���e��W��#��_$��u�7K�ڍR��,[�^�9��ڸ�M�"�����d�����f8���|�C�/}�K��iM)k�q�8���CY��!��d���z-E��8οv��
��2�k���u�����餝�{�	�L;%Z�,��*���M��NS�?N�'c'L�t7��f���߬\��a�0GaM��b.�%%��d���ʈD��i���G?�%˖J��m�/�P�`�_�������X)�A�Y_����΍ՊF9m�4}ˀj��9�ǚ��?������6 h��Y066�T�S&�	]�N�6V�p^&P̪�s��u�]'+�-�4�cY��%���|�;
�P@|n>����o!-}��2u�x�PN^}�F���¡���s��2v�N�t�j9�'ɻO��x�Ң�jo�,ݻ��_O;���/�s3��,���c"��l��$���r���b�G6�4K{{��c%.�iY�n��sY��]v�uO�n?��M��/|��ݢ�������8�8|>�я
-�xX��o�߰�]�~�W<�ޠ������Z �_5�=�/�w����U6KK���c]���'�3�����e�r�#�|U�'��������t�<3q��)��eu��3;Dy��D]M]��Ʉj�G�K6<J2E���g�f�*��?��Mͮ�S�(7��_�y}[�?y&֏��8��;�	 �~XVn[�&\��� 5����8�aj~��9�� ��bV�YF��=7� �?zf��뚀5*�_��<��g�^��Nj,z�(=�Qj�~�U�Ę�@��n^/O>z���,;�N���AW�?&ٌ��Eˤ�v�4��$u���ǯ�V��FIgw�^kŊ�zn~�����h�l�0�k���CW^!�pQV�\*?�k9��äP��VKWW�s��jd��ViZ�IB�zY�z���!�)g&�5�\SZ�,z{8ַ�
��ޟ$R��8�m�9}�`���s>��� V����5�	p�u���o��匇�EI��֑���
:�!
B-f$�k�Da��3����&�}��ɪ�O�?$!AcZ�?�H�\J���7,�bL���;!���_�1 v��%Z�aS[�UE%t����mƀ&b/Ӝ�Й��|�R�P�7��zt������$8z˜�s����\�	�q� �����H;�()s��}[�:�F�"�L�.9�i�t��gȧ>�)u�ҫ��k�U`��K�B��&�h�x��e��k/���J�<r_i�4V����1���l떥˚%-׷KgwV��m�caٴ�EE�.ݲ_���Vf�h(4�=gϖ�\}�Ĵ�C�����;�y���]�~�jimkQ隈�K��NY�z��r1y}M��e߃T�ǼE�n�Q�>X��ӊS���Ik(���g	/��@7�v�cK�qmAT?����\2W��?�}�� JNi����^�+ڡC�������?�q�u��LN<��D�K������|�.��?~��h4RD"�!j�Nϗ��d%$4 ������}����#	��(1��|G�l��5Do�������M��F� �ti@���}�!��1^>?�uW~,�e�o�I����_�m��˵�"0G��6?�o%�IO��í�i�Ҵ}_0r?8|���<��#�<R-�;�C�.]�S��g�(�����<����̖q�G�kK��K��D��saye�r���ٕ�L6,���:=j�tv���C��0&?:�����n���5�5������~L�j*f����ˡ�'�b��Z�B
���i��M����뫤�#/k��ȱǟ��?���8�j4R1G�q�<,6+&�]w�UJ��}����M��^��m?k:R�R�4.��k`rSBAk�����x�C��崺'��2�
�E��ˠ����Z��K��#WKD���f%�k�p�E��M�o��u�d��i��O��JW� ��GjS�;res���Y<9��\l���%-=��C5�'��W_����/k}�����WU��d���b�ͱ�),�}_\������[Pۦ���%
ڒ�ݞ/�K@���S��,��^������Fa��^��P�,��PV���8� �gs�Z����(k��a��iz]:�h�p8"�]=�|�jIeD6o�:\�8���+�_[.w-�/�5�m6���ܹ��L�]]���]�F�{�{������ukVJwOR�6��\�Gyr�$ź��U�o��Y���רs�ŀ���4v��v�J�{�WZ���A{D`��㎅R��s\s�j�O;.��JN Zd,���u�>���xc�����Ւ��q�:)3D�E���u�jA�l6%�t�$�Ih�g�Hj�<xϝҺa�L�� '��Q�O�.�T�GE����{�i���	z5��aL.2Z
�1Z�!-5"�z�<����_��������C���F�;��sh���r���A�<���a�>5����l�}��6����oK>M��K��l�K֭}U2=mZͶe�&���n�hm]��^�$[���ʵr��W�����p�N~��?�/�KF�%����m��8���m��+���ƙTJ�._���$P��d媥�|��QL*,�t��5������3%��V�1swV$?mq�qN�iF�C��x�%n�E�B�s˜J��ETqkT a�泙��:���db�5;1W�=�5�kj��'%�Z7��U��?�u~��-k��1�[�y��w ���F�eR��vK,��!�l����r��ۥ�y�4L/���4��O��H������<���2�4²q�a)(��B�^r�1*z
1	'F�g�)��w�-���Ev�?�����/�}i��Q@��?��X8u�@���9�9���/��ژ�3�����M��A	%�GK8�q���7ȸ���N)Ƥ�'#>�;��?�s��~��ɫJUϠ�b>���cG�YgΓ�;X�]�m��i���7JG[Ri�P!$�h\�L�*���Qv�6K+C"�)��׿�����x8�}48U� � ���4�����kU��*�O��q����Z0*��%�i�OKWG�߸�E����$	�Õd#;���@�/���S��f.��{�w��х|F����%%�L����_�*�Vj�ƹ�d���E���lZ�ZVZ�IT{���/��/���I12Jr�Z�)F%�-�L^�Q��ǷH"�V�v���b���,D��2F��GI�)�����w�h�믿^�=`N��7�B&5��x,,�L�<��S���OHw��E�g����Ւ��s̱�����3V��^�Q_KJ���������++i�tɱH���0I�s�<y�[���DL��Z6o�H��+V�����HmM��7^r���?�L���ø@�RY$h�˖-�Tp�r%j��vq왃W��ΰ��_� s�r��O>Y#���:"�Y�+�fZ|�UWT�z�5�O�1��<�v8���N�����*g�{��I!��P!-�ѼD�ݒ�l��~�lni��;M���q�$�FK���Dj���ϕF8�5��/Z<>�0��:)D�$NH�>��:���R����)��H��ڧ�2�w��ه~�nԜ�D�QR�`�|nV?�d��Ib�߽�ҋe��	l5��sҶy�,Z���\�R�'64(1z�X]�������=��qB>��_��?w����+*�?tN	�pxf���w�q���{�)��u����%� �ߵ�u��IgSZm�����-�>Rn-��+��� "p�P��/�+�A����í����ꩧ
U�Jt�g�����|�s��д,�?��I�=�y}���~*�%�&M��ft�m⡜�r)I�Ҳ�y�!p���S����K��ه��O5h��<��#T �HB��I���ȑmIm�M�em�j O���Ù�ߡ�7[o{p��c>9����M�+�y����^�����l��o�8�!� ��sl6�ў�T�em�_9.��+��������Sa��1�uw�q����46ޔlO^^	���IM����Ak�\CC�w�}�|��%��C(�鲓��K�_��,~���q�\�߉r �k�]w������H j��3����@�[4�j�A�ᆪq.�K��h��VD�B�}�1b���E�S�`�M�X9�� �j�ѨjN�\A{&S<-��Z^
�n���G�R[C7��� U"q���?Q���$��Ȃ���91�XH�X����G&�W�N)�"�R	�X�n��/�},J�֩	�сo��/L @�@����~s}�].��6N�i�2(��f�TAA�US����fy������N�����r��i���8����HX,��.$+���̓�8q��;Fv�4YƎ'�LQZ[��ҲY6on��x��f|FA�h���O>���illT��駟Bİ
 ( �~�����G/m`n�DS����@�NA��k]i�����s�nL���D#��N1��
��pQ��٣ɴh���ҔF����fc�*�e�xI�Y�G4Ɯ>�Ez�F�bk4^��c��3��(��ZKH��[�C��ܕs{i���\@ohhJ5`�*{��k�.�{([w�y���`_�P�~�����t�"�&V�J�n���"��YY�v��X�\�֮�J���Je8�S.���z'�[�gNc�-���%�4�^�ؚ��"�J@K@� +@`��"���ʩZh��l~��Ԇ�BVl�c�.���`IahF�{ktMY7��(����B���-�6���)�ઍ��E1��r���"EpÚ�[Q���h������x�P�P@e!����I|ύ��U*a�`�--����`q�V��O������'�Y��	|�����Lk-�vMS��������5�<[�4i?1��k�߯Y�ܧi�(Y�� ��Z�~�i����I�$w���to�M��?�>�����̿u]3!���YG+\�a���^T_#�g����Ȏ�N^CE��j�P��ҕ9��<@��tJ�o���n&Ο�Ë��;�s4������Jv��	zr�i�Gi����F� ��Z>����| �WH��m���!� %�+p/}��n��p^.z� 	������%V/ޢN|�|�1XL��s~9 ��FeP�pŅ ���=h$��mnݢ"��Kz,�B.�^B΄{�롅㿢�N�����˪�Z9
n5���z�)���u����_�@m�@f��,q�G�PG�:��h�֢p�X������2��:��]�����ޖ�����ی�i��)�
�1���p1@ӌ� �@���O'Q?<|8?٢p�֤�<�[h^��]��Uz ���瀻W�@_-�-^[&ܠǀ+��ZVV��IT�e-�$z_N������c����7��'�O�:a}�R��i���[-״{��
h�\ֵ�t����,b�Y��+_<�ׅ�|���z_`��û���,�J�P[�(W��qƫ 3kz��a1�~��&J�T�=|���A�?�A9�c��K/U@�o�x8A��"G�h�Czq��r0ƔI���}�`D��@i5�Kt�o�M;���(�JZ�3�\sj��X�l(8@�l67�  O��
�ق��P�[]4�7��0���5|[ݴ�ܒ�\��`ӻ�x	���m�KTSp�����?98�X7Dy����~&����5��E�JQ;[�oL)��>��iHBt�����n��Ÿ�H�p��j���:�4�H    IDAT^6�����2�+�5�K�'9�zDd��b��c�ҺY��j�X�{3��"�'d᳧���Ju�Z}.:���#��t�9x�G��6�6Wt��+; ��`�=[�}|�|;��_�K���7.��V`����n'��3Yՙ��d����fZ�{u�Z��>ڲU[��>�?X�zەuc�����7x'h���m�WI�!ʧwc��p��1�w[��J���T^Vc��%�k��_恵u�ŗh�M>���&	���
�Ma�3a@EJ4U�	pn�QiBd@�Fnf������)��oq/�X�:��t����S���1�����o�� 0��>y��'T`�z��h����"�����E�Q{<C+�`֎�OF��C�I/]��:sQy�·o�c�>[������ι9�l��o��  ���X���p �x����X,�.O?�^~��׭ҡ�c@0��g�}s���������ӁƯ1��a�Q��������"��G���;�('�P��pf������b@�o��
��'��¾l��Y�uiA�Cz����}�l ��?�x	p��d��p֟�S�'%��G������W��͌lo��Qg��4wb�*X 4�D�'���R���_�}�����@@���9��}� v@��G���ZtE��� �~���V� ���<��C=u�IL�s&�h�����O����eԉ/ }��Ea�ꄘ�"8,��L��/��m�;�;�T���
4P�Y̹:,:�D��:�0V;�؂�q�����cJ�O4`ͽ����;�*�"
(� �D����o�� �w`���h����?�.��q5˭��ӈ(p�B5RR���&�O82�o �y-'d8�i`��O�:���&*f��U}���n_����e��$�@���k�6�̀�5��B7�۲�}F@��7��+&<��nA�8G��=VYw�y�Sm���f.�&y��O����������MJ�b�3������a��LR�ke!�>�lQ[g�;�/�7���J����~| >�n�(e�z��Q5��¬%��Q�1��s�å�]t�}�o����}I\  ��唺/�pm���������ș���?�����_3A�s�2<�4�<V5λ�/ � D���0�(+NL: ��z���� ����4\	i���V2
�ǜ�|��?���J�H��!��A�x��O�Sy��ϕ�f����5��R	���uNc�k����RþeW
�E����?т������RN�����Bä�.���-�@i��h�ij7�l�:��6�����@S��z���s�/�dN5{�&�M�0��ie�)�f!kV�m8���n������r�>���pL碆�=���%[�J8A�4����0"�BX
9�/$R��L�Dc	�*/mW��_*'���B?{�y��8.?���8����KNK[8�c��I?���eo6�EI� �|��@ͨ�lxr m�g�]�����a�a�s�lH�9�#HL�<;~�_Z\�{!�s�� �K�,�I��Ϲ�[��3Ӳ`�Ͱ�Z�e���s����d7�d�������{F�1ɦ��Щ5��Q����̿c��y��:Zp�ߪ��¤ɓ.Zpׂ;��q�)Ù��w�6�ؖL~�R�'fN"~])ˠK8 �q��a��ٿ�]�͇fO,���k�+������Y�0�!��6��5Sq[��@c6*��}b�)o}Ѹ�t�d#͔%k6�I(z	S3(KW.%�xL��^��6Q�VsQ4�ׂ89��3ʩ�.kkH�rBݜ{�xUt �͒�*<D���^[� �  �Y�+%Rm|>���-j���c�Um0��/~�EȬ*%�t�Ȕ��B�t��̱���Z'�jWe����Y攥�.��Z�|��֪]�,�r��k?��1A\$�]���ح��+	�\М������`�_�F�;����4�JUOJ�(_t%�'D�g�M�2MC��؝"o�����^�|�K^iO�F��c�Μfl2�M�}5���˂�Xk3K�a��U[�&�q���������E1w��VN<���6�̉d;3RK(�Y��$U�H�X��E�%�l��Tid������u�����й���F�VQ�8�m��Tm�������Ǝ[�!��	�4zh �V�U��������)>����D?B��¬v/}}�=��A�;���>��7�!�W�����#6'��Bm|��9Pko[���y�@��+,�#1a�+f�k�� R��y�{�5#�a� $<��%�Y��VUJ5K8Lq�ٜ�(e�WT.F��?gn?��iܑ+�dS����շ�dRZ���C��8P�O���@��8��^xi�����Z�ro���ݚj��y��dr�jf6��a�Y�C9f8�����gt�J!㣥4!~�	0*�����͇%F�|`!+��uP��Ϡ�@��_*�a����p){[D�k���ԓ�V�֦t\ȅ�moڠ�|0a�٬C^�	E�0%b�V�l��O��F#ڇ2$��n����%�O�ܼ)A?����2����]ˌ�,��?^3�V�����h-۷v/%N?k��9�� ��w�]��{�}���N����K{{��{��e��Œͺ^��TֱA�J��

�]4��;�R�:������ɫH���l*źb�Tr�a�hݝ���S+���,6߲	y�񚄴%;d�UkBR[\��mE��/Eܨ���c�ir�J�/	_ֻ��6����K�υ\�����.W�'�L����3Q*#񀟌�Dr���t�R���|1T��C��Sh�oξ��B=K!���&\��;�Nf��R2�ZD� �q ��0����Yw�%��Y�J��+b/+����/9��O��yC��_�B�q�R\�똓�|ù?C��ZG��w(g���N��\�=�9��bn8�	H�S�_���޴��#��|*<���}�q:��	���K�6.�tZ�@&��g��U~�Qio�T�ɯ5������No�^{[�>9�F�Y,JM<!��V�={7�䒋�e`&�a����SO��5�����{�m#���J6_�g�yFc�-ӏ�/��6������A���~�3uH��+����d��@Y$�Ql�u;�SW�P<�j��#����	Eb��B�I��IM� ��aɤ�$^�L!+�X��c����A��6*�AK���� ��j�J �2g\Oڅ�U�AM�f\Tyd=�X�o%��B��k�s��À������Q�?k���,4r�܉'*��7fv/�`ʧ��	&��#)���.�0�����=k�Z3������_��SOy�~�!:T�m�j��e�/��!3f�R*ߘ*�_������haT�LGt�W5��9�Ǝ-��8]<h_�(U(d���<%�$�6l��-�ƍ3Zv���t�2e�n2f�x}0����I����9I�[����EL5)����~�#��6-�8Zs�j%V9x[V�t���|ø�J#�;^K �0��X��ĊiɈ�:����W��nA*v�[e��骍Ȕ�M���[`�tە�_^x�����'K�~�9Wˆ� �-��X�o�X�<C�A�`=0椯z6}]���A�@�ˢָo�Ws.�{�t���1״y��1׼�s-���<�߫��P�����|ǯ����|��=��x�;$��X,$˖.�GDk9%;�5󺶾Nv�<UN>�4�y�LIC�f���C��o������=�h�3w��$�mWW��!T��#�K.�PR�.)�R�ʫ�ŋ$�s�(�X�����1ǟ$3f�f	���A`a�7Z�O<���{D&P��/��7߬ܧ��i�Cs�����W��j�_߸^&�oP��D���D$+�LR��V��rӍ�	e�x��g�#;7�(�Z�,%����JqMV3�W�O�GKw|�d£�yY�k哟��$�W�����b� �8���"�|筽g4���Eq>�j�6&����9�~���ܿE�Yč�*�;��<{��A�ܱPp�c�0�F��Aik*���D%���+�ʋ/>/�������b�����%��%'�����Y�����mwܮרV�b���<`R��!�/�lJ^[�P�lX�$�74�:^�Ԥ!ʆ��;���TH����j�Z��#�<��$��D�G ` ��Oa��ú�DYT���+,΋���b,Յ�^{P��x^_șF��& #�M�0n�\����œ�	�%&]͵J��"�L�����K.OrRX�4ΓS���h�q��_��Co��~U A��B��;�����l^���~�����߮�0+��
~���`�E�Yh�i�vߦ)݈������ޤ������n�F	0�ǀ�w�o�Է��<��E�*{�֬�t���.��Ȕ����L�SR��e�ڕ�a�:Y�����N('�C[7wʆ��RW;V�zϹ2k������������s���P���&7\<"���̝��d��#�45�����U2��F$��_��^����%��U�WH6�rE�����eg���D��w��o;^{��`q4A� �l(6)�>�Na$:B뀈"��"��h�9�q0��Zp�ݶp9����1OY������Z�F5���)��/I�8zIB����N�����&���ߓ\�[�Ѹ�i<K�M�-�|t�௢�^yu��[��u�����L�Fƕ
�1? ߂{�|p�U-�
��=���QHe����{)�}�yM�X����	���P��Ox��vO&�8�w W��r�a@���57Ա�I��snj#A�|�+_ѐU�a��?�����ʻ�<��?�S���'7���>&���$Y�f���V�p.$�tNV,o�H�N6nL�1ǝ('��?���^��%��O�o���Gn'�*�O�B6'{�>[���5��꒮���}�rһ��b�G�4��Q@���I��KV�l�t."�W�ʁ�5�y��8���Э�;���A3@ۇ�4��6���
Vv�8},�e.���ð�B B���{���-�&�T�B�����w�!����$!�?��$V�h�E��n���}�����eΜy�ӌ�%O��W���ުm~7���.+�ՐK! ��=4C���R�4������]E�WP���]�#6e9	�4���O�X�A�'�0���<M�)ꏡ\[5�2aPm��ތ�7�f�0�i���s�Y��y���/jH)�$���sP�xAa��p�z�ed�����
��M��Ϗ�J��wW�0a�,]�DR=���LQ^Z�D��'JSS�4L�.W_�q�������X����-�����G,��vz�w�ے���+�
��n��U�R��>������C%����HGgR%,}f[6%��i��N��h��<T�z J����}�Ta�nB8By�L`u6��f�F��z�D�+Ui�V�Tw�F�u�Y��EW����� ��8d��xp��J��qh?G����-�~�
�jK�b!,�PN��E� �o�����wϝ'Sg�&Y/%~p���f�'�lU�i����[=k����W�������@ɞ�Qp��E +��h�*�O^�L�[��� ߄C�1V^v�rJ���E�ʩ���R�-�g��k�Q9����?�i�+ <�[Ț����<Z_�җ4ʏ}�g�}�҈�y���SO> ��L�0V�-_,�T���;�e��ՒN�ds[��������F�+������?����YC#��46~;ٞ�XE��Y3f�G���$�QiٸV�ӯ����p8%�ׯ��֍J1Dc5���)�[$����u�2}�n��O~R��L�u�]��ll&�Y͛7O31�������$n�\�b2��-�8�*��9v���{�:�D�X�����X% ���u���)�>+�ʲ(Gq�Z?�A1.���
�;Ϳ��N������Zy��g�ԝgI��;C��5���6�}���F�G��>������9 �hno����`�?XW<����)|+�5j����JM4Z���T�P��}��0�V( v���j�;������w�Y��'��	�TA�Pv��i4�F�S���6�oʔ)�-W�Z"���>��ݥa�hy}�2I�;u.�+J1&���H�^��9�������_�DM��(��?�ח/���✹s��L��/�W���ҢL���|���H<�h8/�T>ho)�es[����ꦉ��=���5�d��Y��SNx�)2w�\��l����'[l$�8�I���eQ���� �-����Dk��PIh$�;��R!�l�тF�M�O}J��7�������DC���v���$�����rىb���-7h=�p�^N��?���:�������k���Y���n!����X5�j�3�ʱh�PD���|�V5�&��	�ٳg��F4~˲-�N�Ž�ڻ��HM�����)(6vߧ�y�{&��V���*�p� >N_,gzPn��n�����3��g?��ww��SO�Fv�e�����U����Q'.AX�.	�H��69���e�Y�HM]��Q�z�J���y2�gräK�ϟ[���__ح����E]S'����-��!5�<���2vLTZ77K&ө��<�I��d�Ƥ�i�,m���+�Y4���n����o����6.)�d�ZV�ղ)����%nX�E�P�j�x��<����(��s^Uƅ	K�x�.��LP��f��a)�sr�)'No���OL�@$=��&�)��o�;o�A����i�g���H�8�Ԟr��^j����4���L��1�޴ȵ�u���/�Ɂ8�yA#P�� �4?+�փ k�5J^
�4� �|fl����~&�����m�������Z�q�o̲���e��ђ�X4��_���g��ǔ��N��%��l�[6�4���O�|(!�6u���kecK����d��p$"x�O�8��t4A�����_����k�q�G�|@ҩN	�Ҳb�bY۴LB����0ц��	��²is�L�eO9������Z�������i�?� ���E��ԤZ6<����M��$y�:O�R_W���7F��DB�r���fiK[�R�Ԍ��lA�����P$�)鍧�K��;S�uǥ�3R���-���;�'�ߩ3f�_2�i��6C�M��<���8uU�7���c�'���"�L���:媫�ڂK�@8�s�_t�E�\�SM3C�T�4p��N@���~�ܔTF�	�ZQ�G��xs����(<p?|�����%|Yة��T�d��l�{����\z?� 7���ɼZ$�|�C���l��j> ��;���
�Y��"�Բ^
���ջ�n�V
��,[�$;M�.�x�I"r�P�k�dR����'Mn�l�]~2�4�j_�,��y���������)�\V�z���<)���	B"�e�<i���]�!���S�5�
����o~�	o���_ %z��g��X���e�Z�5�bc���J��U�I	'�?�X����
�!g*����"!���:[�q%a��J�q�����~����K/���~�kFr����3.��?�W-�j�<��s���*9LK*����os(k�ݾz����o��,[[*��GT��M�lx�>?4dӢx>P`���_�܁�P�cn�u�*`�Z������`%� 0��iԈj>`e̕�c@��8��s�OV =�q^�!�,ɑ��mfB��"֞�� 2V+��t�2hå}l̾���p/���P����?�Q8�n?߳,`��L��1}����Xs+�.�t�GǬ�%^#uu�d�]��#ߪt���O���n��]�j�W���{�����2|��O�E�`�Q�	چ����>��j�(6���n�g8>���+��( �w���i�(����v�M���ok� �C�fX3�j�OooY�h{i��U1/�HDk�G�Š-ڹ�x)��AP����+�B�h��$H�
V��z��,ި�%���K�mG�Ux@��Mڹ�y��k��Dr�r�-�ӌ騂��2}癚<d���9T����0�PL��'>��>	hWW	.��-
�����@��>p�* �mp��    IDATk��&���7��u��h��#���/V��^Z�p����~��G�g����̾"J��s<[ȭ�B�%�k���?�#t�$S.^�Z)+8̧�|�߄)
������gF�|?sl�c|�#�Ep��1��fT	&��a��B�{3G=Y��~�3�j�ܴ����~�z�Eۣ��+��$��3�h����c,^k�d�Z��駟��k��4���� ���4 "X�x��u��jR��BAM�bT˰����G��Z$�m��R@A-�E������\Ahd?�O���_*Gu�V��������z���yN��M��p�$�����&��j/_�g-SX�4,M�"������ |��!��ZrbEdQo��Z�L������7ARm��ל��@?�1��/|A��=L('����� <��K��I�:Q#,��s��!b���D����b>+��wh�}�@����\rnY�����!���uڃD�g�P���<�W���=�����X�p�V���������ϗL^�\��ˊ�tP��zݖk��|Nj�Q-���~�.�K#-�)��`�B8T�����2��U�����S��4���4�7;�w�v��ш�� ��'N{SK�
�lp� �� �X��}H�k�������v��m|f��� �;��wܡֵ�a�<����r�[,,�
͟(����O5�`��Y����f��v��V<�=> � ZWR�Ǭ�� ��������:JKD�]�|�w��P�
�C��a���Ϳ�#���1�����2��Ĳ�X��e�Y�"�3�m��u�^ܯ�c��]q��p���,�j�8�~40�3�@,�El�j������6ܾ�����I����4&?Wt�xE��=�?�գ��}�A���ϣb�?��(�(�or����F�F�� ��@��}~�NZ4UA��������?c6�Ф��*Y�80�o�k�kXn��?B��g�ؗP��?`Z�6��傈�s�'؀�H����&�/��BIq�Z|�%`]�u�����1c�j���B�h>~���a�U:ۻ��������t�Ι;����k'��Y�.6̀��$eaqF�w��O:7���/	���-|�-��P�;X��@�-���>�C�@؄
p�QI�H�����.4w^�܄�����4�j௙����>�8G�>�������i4Ž��{�/�9|����g�h������_\��v��m|�4���t�w*M⃿s�;%��
6͟=�%C�ǣ�C���?�����/ �|&��M���m("�Ц��1v�V� ʤzJIZji�M���ʭ����b)�7�2*��N^#4ο��d{�r���s�ol��i&��AZ9�ɷ0N��i<��o��,�dq�!��ބ["�z���y���8���P�װ[l��4���?�q�h���p�M���������5ZY�h����\+� J�2��?������Qee�.��(h�O�~}Я�����?��1m�/���"�������1`6��2>ބ�Y�������-�������7�Z^6V�5�r�+ױ����ƹ�?jK&/��&�m���<��o��k����w{�v<��Y��%qY�-t~�>�[A��Q��ĩ�B�9�q�.^���M�/Pp_U���}x�,h��q����ڧ+:]��1�o���i�����RS|MD���$�ֈk�u���LR"���3Գ��7�Ǣ}��њɏA��e��r��ڱQ2P��	U���t�6����iS�6�xߺ�Y�$���ri�����m���9�y�ʼ���{�
V�k��_a�̝ss2�~i%�f�BA�0p�T�຦hT���^��_mCb�
̴R]_/y"��!J��x��L��X\2��d�"�0�D�.@�8�[A������ΔS�}���E�@���h��>��{6.n��z��WK(H�y#���'Ml����`��U+��'#�N��f���LHl���3��k��i5�xȤ����󀳼����m�vaw�]��A��A��A4R���&Acbc��I�Q�`��&%	b����ԥ���l�;;����{��s睻s�.;�J��������k�-�9�9Ϳ����!%�kF}�9>�|QHϿj޼�_�I�%����Fm��%�5á�N�ܔ�ɿ}S�?��6fa)Z@בE�@�,I(Q��H��Gs:�cZO�h�,喖���%ʫP*Z�R5�������Th6]��+������V�v�ε���\�/9|�}F@�n���M�(�v��~}Y�M4�a��Z��V��h� �Ƭ�F��|�
���袋<�h;!��C��j+�o&|xV�}h���F�����^� ��x�o4WR:]	{�4ք�s���;�����O@��Xf7��ȹ���6u�5����%�R�m&uX�Z�l.8�� ��p���eZ[lm�z��h�j��?_1�?�2�P�bs:ϱ����8|Pr��ܣ}����O�������<շ��� �������LE7L�?�>ǏF���u���B��{z�����%�ܾLʎ7��	%��Q\X����FC���9��������8�I��;z�	�����J>�s�x��~��i#��8�CŞ���yS�X���T�/4�UOq�\R��l%��$y�����Z�>K�zp	���A��������ߠue|�AAP��R�j�~S'�%��t�3\�
ȎMm�;֚���v `b��5Η�#�#��N4��*�������3.J��b�wliku�u��Ͽ���xĴ�"���hA�s9�3Np���|���M����#m&6�M@<�����,�ac�h�x�����-����I�!L5�#��*��[X5���+Y�J�}�m�����3�i�Bۉ3�8��r�EV��]�_p���C=�?�Xdn���_�MH�(�E��P�f/�'M>�jDT�X׏�n�{������Xo�C����
��cy�0�^�Sۭ�lh���'2��9��4��E���/�����V�o0��t��5{����ҠK�ġV��q���P~G��b�+�k<�(MχD9Gswm-�,^"�Z��ʹ�{6��įJ!�����]��L.���J�5��H�/UҞLv�)'�e�����3�-�"�'����"�������6���o�Ǎ�}���B�KȺ���M]��KqX*����v��I�Xv�B�u�l:���0�XWZ�)�c/�J���8��ⱎq=�SO�	W�Y6h����x���� "���O�6X�B�|5m���D9(�wSP3��뵃^�*;������L	��=ے��׮��]���߽���x�0k�h�T�|�	�ٕW\��>p�.<��q|yv#Գ��R��/�'��M/���2��V|~�p�1�"�?�"cZAʋK�/�����h�$�G�c�����5ݍ�JH`�C2}ϦS��M}�?�y����4��1���=��Ϝ5���o�����O���Ku��\RB�0;@����o�Cʈ���`1�/n4|
�Qȉ�Ʉ�@M@f<�F�?ׄ�)��v��ϲ9�����Vs�fq�fF���Yw�z�����z��{�����Y{�X�O�y��!;��W�UW_bϳِ!\-ZKe����J��s���iU���W�3�c���t.�B�� @A󧄂�q�#s�5������(�&;X��W_I֬(�p�\@�84�,��]2ӳ#l�7�c#�����*����>��@��G-�O�'l�$�������R0�s-�P	<�/`
�#h�0�ͪzVK3g�x���fq��c[[��f"r�
���a�v�y��C\���t�Ig�t3�����͛�l��LUi4 ��>�!|�{��@�j(e]��ߴ������F��JR<�1{�l���7y�>ז���j���3\qՕV*��b�h��p��d�z����r�Q���5=`�r��U�[� �f���v�yo+��V�T����A��0���Wӓm�u��KLOp�ui���5�`�j ��8�\o������̈�\2�4V��I<�l�/�3~��j��b ����<C��#A*��`�
��8��C<�u��h�D�� �)W��#���O<a+W-�r�j-�4�
ax)��G�q�-�jub����}���/*;Sj����zՁ6iR{�$
�ļ�y��/U���@���뮻|�dV�V5o�6<1�h&D� �|��ޡ�?	;���aƳ�Y���Ѵ��n�lB���>��������L��'���כZ ��
Dۭ\��L��J]I3�U�͛>����L�ٝ�ێ����?�a��L���nV�NVP�����~�%�U�g���0vZ߱,v�}�9}6ָ`�r�r���Z����EK�BG&�;{��9^�eŚ��R�8��c^k��q��M�p�Jh���6))8���k�y������B�`��ϴf�ђ,�$`+�'+fvg���=�kE�Դ�JH��q���/����5�b�`}��}r����͜i�����=�2hȿ��/] h�0�u@���c�Q����3�\��뼪'�%,b����Q����k"ph�'�P59�c-��P��Ѿ!�����nSuJ�ͪ�3+�Ղ��^Ye�b�}�Ϲ� M_�ﶓ+#�[�ol	lP�2#�9�����VjٶֿVB�
�$����,�3A."-?��a/J�b��aQd��5>�	篨(�Y�V6�����7	%�1�|	�gǲ+�{Q���9ԭ 1��׼�Zr���������f*c����,C:CK؜�E��O��Z�iߘ����Z�К�9�v~��;}#��}@�6�LV����㏵r�`��m����k��8y�n!���v�񯱝v��
�Р�ʄt��s]��G��u�8���?{�w1��5���as���FĢa'�X8��gu���6�O��]v�e��?Z�g�j�b�r�\��]�Q^e����͟�J���?{ι��n������V��ץIR�: ����.Vi��c.m�1�����V�t!.�\�k]+XB R�&i��˾�}�q(n������jo� ;�}O�q�o\L�Y4�>�o|�y�˦-C~M~�=�Я�_�<�T��ε�Ge��q��N/R���ݾs˷���V�X�q����z��74�R1^��:�����k��bi�2���X��~�z���V����S��p¤�מj��� ������pg0��'�OO,�R�Y 4p�q�<���G�g��g<�����(�+L	�s��$��IH��ў��
GWlֶ�ؿ|���:"O�5W�\����W��o�w�� �v;g��t�s�5���9�T{F�y�����
�l\�5���㙻?�s�*�k��M�Ԍ^ �Ϛ�?���8� @q,���ԱT����:�q��g����}�����}�q�{��l�vKW
�j�2{�
�5����!�r��'Y��SՌ���cg���aͲe��%	���	�1s�w�z�����O>ڧ�����ο��gҡ�+���;���-�.��yOY_��\�Ժ׮��g@�kw�Zg��e,d�]7��;�Y���ַ�A���B�w��S,, �9?��3������cNqS.�)KRB��#�,q�Ҷ8g��CSH�,�m�N����-�	!��R�Z�U�V{-W\g����߸���m�s:q������sd�R2�[Ç�s�HX͍��
�l���_A_������l ���j���O���O�aq7����D8Wt���P����3��~�;q�����?ֱ�p��ҬH��"�d*W���Ъ�O�V�(����~�"5g�;�Ӭ4�o�}kl�����m��.�e�����T���ݽ�v]���~v������6�c�}�;߱_����'�
�fw��9�����!��������v���K=�e*vם��1Gf}�����g\��j�[�.o,���ڲU�v��'�\��ˤ# ���ڦ�zϸ�hw�Ue�}��x�����{*�&֬�����X>��a�Z�)�-�O��uLF[Iy��ʖ�>˖�Y[e�Yq�}���Y���X���l����
�i���Ӹ�뱗�~�ӱ��Ib�{�i~R�:d>�V�}zZ��W>~2>���W��ǳ�F��Haoq��gu���-$���4z
�3�{�����k�j����7�[�����i`�_|ћ��4�a���3�K�=kJ%,xƏ�㾮��2��㿴�P�͜��=;�i[���{�
u��E�ʴ٪�n;�����ϲt��~��Cv�w��@o���hkuBk��tv�SOO�Ɔ�5��*��]��k�=����k��w�f�q���Ru�E�\_\���A[�d��*��pq����������Gc����8X,��;��}�+�WZ8���ŋ�O�bO��9�6u��<E+(tT��4�X+��Q�f �3,��ђ���Gl��휳��JѲ�!K�z����T�Ǿv���S� ��Yi��W�~ɴO<P�ų�ʈiJM������g��d�>���[���O�����'��-�y�3oФ
z�#��z�OIg8t-��3Xԛ#�^�Bk��b��
�_vɥ����}v����4�~��&��k�-�6Qqt\�b�=���۾��bS�L�矟�ډS�ٜ��y�b-ֽv�v�y��򫭭}�[7}�f[�d�V�o�@fϙ���|��������o�\{��Re[�����e��z��}�յ��z{���U����]��?X�EK��+�;������c�|����BF+�ē�'��{�mT6��O⋇��vl4��Q��{���U��P>�=e�4����Wmr[���!K��<�kš>+�)��\K��������v�G$6BbD�n ��,0��|b�Xf�+�v���RSt��h�/��'��3k��o}�7>G�˗��%�?~�����X�ƲҮ��Z;��|�1o����󛥜�����I��}��uk�zT�BTIY�?��}��i�@��g���{�q{��w��G�	��>���Z���Y�X��O����|�������g���]0|��_��_������HMh���9��?��������Nv�uW��t������)'g�L��?����>�����l��%V�v{qI���+݁��ô}���_Kؒ�/���ooG}��s�9�Ezǝ�s�@5��&����n���8&�%�9kC��p�'�(sV��j��բѰڥJx[&kE���]3�y�b��h����I9d#Rd8HkDZ�f7}9O���F&I:��Yk�e�6z4��6�XJ��v�o�.�x�Y�H��͟��3�я~�Aozӛ�W�j�*��>�яz����>����m��=��o큟�eG~�M���-\�B�0��
Q:�b�>���E��)�G>�	�2y�����׾�5���s#譭����sf$����F�O 6k�v����`�-4#)��}ێz��V�5kWY��5.$hX�b�J�^���dE�q䱮ɠ�,\��#~Xtj�ƽ�T� |��g?���{｡v~�����?��c��@�r�nC���%� �8�˰��L��28d9��V��{���� ��A���}�a���w �7��J���d}lrix<�k`ԉ���l#P�(X�P5dU�Ҋ�c�?~z���������� �F�O�s�y��Y�{���_��g��P�(r�]v�;�|?�����O�����U���w��{�lmm-�l����'!�<b�Z���t��s�}�ʫ��z����^�%'�JK��Ϛ1���n��k���'��L�omi���n����暫l�=w7��#�����Qجh]���W�T,�C<��s�z]��YW���~�����;�?��O4��tLS�s��n���������8�R�c�m�m�Qj����Kg���њ��gCW,GR�ӡcX1]���,%�	�䟁2���ޗ0H�x���@'p�c��lL��
(    IDAT�?�K��(IP58}��f���۴i��+�� �i�8^g��e
�D��p�^~�e��>��5�>�����C=�� �����<��`�|������ͯ���cOe=�z��d�
�Z���/��?�Ֆ˶;�t��_�tv��CMY*�<s֌+o����N@����ϤP��M�o��k��%m��?c^��&Y�R�����1�%˺l�=��#�<�@L0Q"�/���F �����O��a2zz�{�v���/Lڗ��I�Q^>!d�V�+��P�V
OQ�7�T&e�T�J��-�.g=s��?)�7raK�'{m�[�v/�:�B]% ������Fxr��(�F��;��ֈ�C�� �G�����-���W�"<�M������W�}~G��-Ͼ�� ����:�i����V�E�����˭l%k�d������)7c��csm�=��O>Ͳ�V��l��η=wH�ӈ�JJ:_uǭ�~e��ء�$y)
I~������ra�Vu-��}�y���?�×�a3��̘1�Nx͉����y�;��mh�Lc���=���k5u�5�M����s��Ga�,.%em�8�-��]8UCMO���:�4 w�d���0%����2�!]	UC�-���U��� Ц`3�x%��Y�>�^����7�w���h�?�n�Z9
�e������{�5׸U���8�������> w�ֶӦ{�t
5����ş�/��gS�~A��;ﴃeR%[��E����l� �@w���[�~�Pr%e���n��ez�m��Lo+:w�\��׿�B�YT�����O�{��n��KG��BU�C>8Ak�Y{G�
�6�3������h��Z<�v�a'g�;&Mqg��������}4�~����JO� m�����;(����3�BMSZ�c�+N�x�>���f�j�rմe�L�R�lE��+�%}z��L�J�@-\tʇۖ�!Z��X����q|�?�S��ڐ��8|�͛WK��8�4���]w��0_(\�3ڇ{�\[;����+.�k�X���G�M��߃F����[
����>$�N�h�\.c˖,�����}�����w�o�Wڱ�g��S���6~�B͠�R3Z�B�����n��扨�&��~g#�'��5�J��\��:�.��"kk%��6���`)0�CC�E��~�Y������MQ�C3!i���������'�͉G�$i�\��@ �s����e�� ;��sN��g��-!]8`d��cx<�f�kc��|��˄0OYX�ކ-��Sx<�����7Y+q�'mN�$И�Q��Q��X��v��w�Ã)ثh�(a8|k�S�u�a�0c�������l�#��Ѓ���q��5�чɞ'a��5�F��cO>�d;�3\9t�X.c==y���m7é�.ϱ��ߙ|#��p�w�(����5���sN����w4mve��7���W��N?�4�o�}|�x�\��0���g?�(����9*�8d�}�;���w�B�D� B��n�{đ�+��	5�N��6!B"u���8�{�>��zp��h�bn��]�A�(�{0�C�q�x���E��C5��y��������|�=
�9߬m�c�B4U(�~��b�ࠏ?�S�[�M���:1YS�t�]p��3N����˗���w�=����/ae��^�����l~�����ӿ̐�s@d@�f�{5ΤP$Q=$xQ�
�5a�� PQ�
�i���%��jqL��S�AN�Ϣ��f���f%��d&�Ae��H	#������R3��I�fB��_��q���7�x�GQ'\?���ˎ;�8��ǧ>�)�&eQ(���I���j�����{͝�WX7�^������K��i��B6��c�?�9��W�P"XZ&?E�H�H�h�7��?�X|�T��k�w�fD��b%�ȐEA��T%�ap���KfS'O���V(B���ڵ���z8w|�����w�?�������0gP:�~�pSwE��3X��@�?ɠ;�s�?ȸ`Q<�����\����, dBs��s:�Н�_Ӑ�I��2�Z�L�6�IP�1���D�9L��E��R������{,�!�����D;xꩧ�+$���U�g3��lsn�|ˎ�4j6�ֈX'�
bwGwRwF�z�IO-�=��r��H�DY:^חe����P�?�u��x�Մ/��!*����N���1|�����M|(� �Bӥ\k�gl�L/��a��R���P��U6�����w� ���W���܅	<K=hk�@�ȳ�?��FB: c�τ��sf���K�O����1���dVk3q\\S�8h8C�I��\ t&�s9����`
@����4:i�ٜ[�ݲ#�<K��Se�e����ޱ&)������� i��ט=�u�{�4O�?���xF���El��'�7 �Eϥ����R);�f�I
�Rb�^�ʞ� 䂕��A\K�B��<#�f��c��N^P?�>��k�P8��b:NV"��t����*�^o�qo	�۪���zgwv�G�'U#�_�Y�˱V���:���L���f�5_���ٛ��f�����X0�zg�y�Kw"pTq�"�bw<�s�[vb͌y��-��ZІw帎��i�zz��@����k��aL�H`p=S���@?J�ñ��艐 H<�8�`�q�(:=��%z�����e�och���I��TEb�h���/A���~'YiB̕�Z��,v�B�� ᭆJ� ����@�q�-��c�T����9�������|��F��+��A����8�J����-���\p����U��9oٲeN� �!�.Ƶ)���q�18�ڪ��,�X��Ġ\oQp��W�Xv-7)A�/kU��h��2؎k����^8S�����?9��e�d, ���N2Syf(�M3�SVl���%tmů����E#�ߟY���3�z�į"!.a,� ?��\����%@�@�1�<�����K44�+bc��j�R�5c�U4�s�����+�����$ˤ�yZ��Fc��i9G|?�7�o 2��<��^d�����Ƶ����t�s���L��?~js�4O=
�+������
����c7��c�����$\{C͸�Wq@��_�[5�O@[��="K�-�t.�P
NU*߃�	n���H�}�e�fp'�[a(���A�j�["��'��MLw���O�_�g�/xA��V�ϱ~�Jh�M�=�;��'�{�ܱf�9k�շ�r�M������9��Λ{��7�Xï�~bs-6W� P���4����z�������2�!��Ŝ�Kۖ[��C��@JA#��M�	L�f���a�|�$J� 䑲�7�.��2�Kg(^�=���@��R&��c�C��P*�|3k�3�y."Ɉ�"�&�l�X)�G�Z����˂�r�eE�;�b���.1:�g2D�T��	�-������U�����������a�$�Q&�%uJ��p�4w)�RP
�R*bZQX bc�Z�VgΚqՄ��sf%�﹬����I�b�I+��%�%�X�/�q}���LҖ:FZ�6�ứ��� ��5�`��e�b�S$[j�{]�Q��1H�;�����k�}��k�����o�|�����p�KQ2^ԣ�40׺�K줓Nr ���?�$3�9AԒ�o��,$� ��K/�ԭ	���.S$���p}�x�l��WG_�E��T YB�d.��2XE��Z=z�(DT�0#�.Z����fB^����ɐ�V�G�Y��=�St�ش�x׎Ώ�0�;j%D86���SF7	�f�w+������6��ɒi%@�F�F҄���8@ I��uo��ב	-gd�o��&�Hi2����^��I0ΓbPԥb�/��͌��o��o\;�j+N~4�v��������!�4.�2 ���_���[n���Ϗ���	'��?�>��>H� u���E� ���p�O�k�B%YƙZ7�?k�+�&�LLKĜ����α�pl�O{q?��P�)����$�>]�L���P��l]W�RI�j���V"O �V[���L����������>�q.�D�
ԳC� ��19��=�QH���o�1標���My�c�&K��)��n�$��H���Ц_AIk,8q�rR�f)��j�~��Ό�ų�ŕ�"��b�������B���ȣ���[G�Gk�}>'A�"f�iA�@Fc���/�Ў?�x��hŃ@��T傡���}��j�r@�0�\�gĪ �\�k�h掁�@�� �i��Z�B�2�����
1�N}��A��k�b�\R�����O�aKD*�%$ejs9B�O[K��9�J�leچf�ҫ�}(�b8�w��>7e=�t����E!庶�:�M��Jоe�H�7��'��ߌ�g�\�M)�C1�|�{r�2��M6�&De���MY4�����G3�5Y:��M��^Z���2XEn�`���_�4�XS��>����$���_�����������?� ^P6��������~F��: ��H�BB|�_p����x�8�K"!��x!<�}xA3Q�W~$i�γG�/��WrO��O �Bk�H 8��K�-Yh��͍Rj43��y����'0K!n�+�)�y��J�`�,��RVJ����)���Vk�%m���-�
���rnsC�s���hj�Y�(D��f�'�\&`a��Λ�=��7���1��] /
��/N��z �OR\[�!phf�5���~΂���#-8������^,t M\&�g�ӟ�4l����e�������C�w�ԃ�'�ZOh�O>������
��K�U���hd�}������՟�ٟ�` �n?�n�kB��~���=a�5�r��w������G<;U.���K�q�G��1���=��8���m��b���L�c!�fU�y��UI�80���2N	��%�[�q��L%k-�i+W
V�!KUKVv�?g�
I ��M��$�������]{�uȍDM)@@J�h�P�"D
���w�ڷ͒�"���?g�PO9[Ўpx[�qlB"7(� x��is0DV��c#��2ɘ�\�SE��h��=�G�}��~#���黥5YL�hƸP헱!����g,�k�Y���a��)����:��g� ܧ�z��J�_�0������q,V�b_�tVׄʁRB�#נ�V�@2�9�nR�@<� E�i��\-���W���شO=�C�S>p�Y|���U�k�Vm��w�=����V�B�bm�f��Y;%*I�*K�:�g��a�w(/���=g]��XO����2��;d�y�1+.�D  8?q��2va��M�3�q�C���O�	�GYh���~�8�B���0���L��Ϙ9�	�̥Y��(&II4H_6ٹ�ז� Px�����pP��<��.���¡x�E�L#8�-�x˄	�F���_^�/�;�28cΟ���
\��g�6�r�\1��5'�Ua3�����%*ǠBݯT� ��b�E5ȹ����|�r*� �i���7���Z�f�U���Z��O;��8�Dˤ����Ҷ�������3@\�;��mP'h�:q�А�,S����u����ڊ]�կ�j]+��Zmw�'§�D�T�X����Ж����c�r	氖���'�x�+�̹B`����Q؍a(��1}�hMh�oV�G`��
��s�:�N8�P��2���n�ZK���|�,��utLu��{���2��Ln3�̖>���駟��R, w��WOc�_�U�P��Sc/�L �����e,�{�t��
�Sē@_}�.�Q\��=�� 8K��zNC&�8BD��d�i�şK�������_�Z�c[��5�nf2U˦�V.��i'c�{�IV*�[*M�i�Ǟ���@��5�O��Rٜ�R-6T*�50�+�T�h�){��Y��+�h����k��?��m�]��J�^�)�9��4�VHyd�Lr<�p�y	N�W��?����;��k�S�T�U�,m�&4�7��$��*!��s;��o��P�![�b�����قE�\.��D�;��C�SN���lk�v�B��tcΎM$�_�_ٿ΅��A��sbPP�q3���P>g�vz��{�s���|�Z�W��}B��?�K
@����]*�������6�4j�6'?���:�F/͚��lTzAsͺ��(�4u�g���/����@kF��^ti���(�_�g$� A"Kgx�|=#�'h��n �{���٩'m�j?�>���l�v���<CJ�t��Z�m��1�Z�H-�ݷ��Y�n��"�m��Gm�o��RC�*g���h���w,ߛ���Z��=���J���-Mt���[�i�C��d���Bi��j�+�B����ʷ_a���a��y��.��ϡ�at����;V`�����#�w�Cה�P��'4�7��_�(��g߽�?��&Mn��U�����Gg��5�kQ1LJ�[�v��Î��:�'��&�0>%6q<�t��ALv'-��@m&mQ��EM!d����أ'�V:p�4,�x����	��T��c	2�
���" �!�/@�˺�8]WB�ϤM*�?��ba�k5��e��Z��H8�&�6���&`��1#��!�3�ϡ�U���~�s�k�ԓ^m�r�����mmڶ;��`ي��M���e�mV,T����1c�M������P���gh͵Y��gK�κ�.�j��ҩ�u��ؗo����X�rV&��7��g���X�g<'�G�[Y� �A�-`]��>�(��u�㼟5c;kɘ�p|rr�Z���Ckٌm��L{͉����z�C_p��9Y��Yi�����|���F�>���ʦ�6{��v�i����=��k���^m^x�z{{<b�D��F*e�Ww���C6u���_��ӎ	��~DgP���#D���	Ĺ��o~�I8����I�
����ϕ���S+������|ST�P��w�ѵ��w��a`�������@1S8fY��.Y /�'*�*�����
J�=�/��"
(~6	.�d�����xw���NT��e3��}�k����J��*Ռ��v�Y;�DҥlҤ)�΄օ8|{{��\�����v�P �{lh�ZrE�Z1���4�c)k��]f7}�[��b�T�U2P��T! 4t��=6��Y/�5�
�V^���}���3J�J�s�8�^RV���.[��{�鹶�7�t�?T,��@�֮[o�춧�~���ʹm=��[o�x XF�O'y��}b�z6�͔I���iӷ��2���w�=��+v�R��-z��}\S��ށA�Z�e�r�-�׽�ӳ5�8���-��ވ� �����pCy�������/x���!�|,ir,����j�c���Oc.���{hl>i��$��<v�BH���c*�O�P�S�0�"�!v��z�N��K� �yLO�7�*�/��{Z���;#g�$�3���<�4E�o�R�>{����I�=���>�fZ�c�^��nX[K��������R��P���´��&O�/�io)YO�E��/5+�[&�f+��K7�a��a��"�ԁ��y�u�A	c\Q���%������2��>����m�f�>�kKY�e�[�x�w9�500d�m�mɒ����V�Yo�\v�t�V,V����[n���h���&4�7��K�1lםw������X�w3�?�y����c\SX�|�5Pu�?���/\l}�f�W��~�b�z׻  z���Hh�LL6� �٘�9��u�U�\킀�!�nEn����8uƂ���?6�v��f�c�޹��6�w�99J�Ҧ 8�x��f��`9�b�&���u�����t��9c���Ɗ�QB1m#��A4�^]�T+���X�H�q�;�3�v�%{%Zt-����
���N������'a�r�U���.Gٔmw���oZ��B�J���th(OC����X�0��{��Y����׻�o�d+���7�ak֕\�SF�	�    IDAT�����_�>ߓg`�E0�\�`�PY�ˏ�dt3�(x0X�KϷ_?��}�����Y��s�u�;x��l�=�س��vؚ�}�������v�k�+W��<�ŋzm��"�W���s���lOw��F���Z.�>{�e�|�u�Mm�������c�y�ў��l�"����	�d�֓�%K�Y��j������~�����v !�����y����L����H<�y��>��x�v0�C�9��scC��[��r�4"J�F��{��>��̝�hb*@�W�t2_
	i�Ҩ9^��|��/��:�,��U��}E=��~=��Gk��R%(�N��_^1=U�p+%IЮ��Y �h�T�:�9�N<�(�z�Tm�=�:�Z�gY��/:��	`$w��������� ��YOOޓq�����Ֆ�-�j���{�k߸��v��b��MLmE�RԍVI<���d=u�Q��o��6/����C^y�^}�}��f�n%�Ս"8�����_�mGq�M�:ٞa��*EwDS�(��g/.Xj��$[ݵ�֬�O��=J�ZM���{���|<�-�a%`��o������c{���X.]�%K_�_��#;����R�ŋ�@G�˶8߿h���ڳ/���~�Wgd�����?\�h��ꪫ<��+�q~��pΟ"]J�  �(�J�l���q�V��ǠG4�Nr��$��o�� �l$H�o,�w�e����˚a��S�� ]O���|�)��m��@�?q�|VuZ��)�ɲ��� _����	�RB���[b!��#�w���W!�
��5�,U7�v��N�לp��J�VI����l��if���0�=X�sV����RgK�����2x����P/��
C�V�H\%m˖���[�ۖ-ﮁ����o�F�����b���_�c��O~��W�r8�x���|�#���z �������~�=;�l���J�h�\������-���Yת^�d��>�i++V)��ӟ��-\�|�*���X9���\�p�V1C�Y3���|��V)z&�7�q�w����UK�o}o����D^�p��*-�pi�~�1^G�����(�t��l6x`�Wac����Ss�=6��Hӓ8h۪�7����? ��;@2wp�l�_��מm)�Z!���UV��b����/�ιd��X����,rBD������B8��X��Q X[��v�\��ƽ�YOj��#Z��F����G���R��R�;o�T�,�1�Q��]��l������9�
C��ɶ۔�{Y*=9������\�t�ޝ���{�X9+���0���a�������
�P�ǭ��B��5��ׇ�|Ya����{��w�XSO	
������^W��f�c��"�W�Xh���ǎ�Î3l��'j��Ht˶�ܧ�Y�J��m��N�go�¦M�i]]��N^�腭��h
�L�J��I�f�d��Km��w��\������Ͼ{�`��]���4����x�R��Zo��%{Ӆou�`C0�ԭQ�8����cs:/�¹3��h��).��7��V�o��f�% H7��T�C=T�×FkYr�rGE�����
@0 ZD�!���zj�E`��gb>w�K�)�A�?k�{B'��  ��L���r"J@�kp�]w���p-��~yQ/�u�f+�(4{ u�_JX������W*���%����jf��b���#Z����ed)���@��U���r[�R��[*I����c�D�� 0N15w�Eفh�W嵳P ?����R���B́�&��ŖIlĽk�&������18:�l��նx�*��ڜ�7�QGo�t��>���緿S��}��U=u�J�&��3O�׿�4*���}���l�e���L*k�\���Zg+��m���|��j-����"�ŵN9���j��{�q��a�c�N��x��s����#(-Sa�lZJ{ �R!�����<�N�����bߍ��f��W	��:�ی ��Z9�ro9��q��g���# }��|�߬)�G�>פ�3k�sE��i+�D�EMd\�H��C�C�1]�G�����p�|�G+/�<>�R��M����J���H����B�E%�s ��f�3BI��uPM	�I"��$y�9GFio��G�n���<R�A@q����q�E�\��o�r+��.�[e�kW���-זAY�5k�=}�1y���^o]��-��oo~�%�݌�\J��w|�~����5Дc���������[�\�?�r������9�_����6�×����O�`���ˎv��o��ӦX�2d��=��Þ���i���l۩����w��;ʆ
%��@3d�C�F0��DBew٤�+N��墕�!���G����?����3��(hȊ�Q��;�K\U1���#iD1���hq��@������ơ m�K���h��%A=)	`�U�
�qM�����x�y���`�p" ��{�zR���� �zQ#	3W�+������'Y���ݳ5*��y�н�
hᐸ݆'
�L% �?k�U:C�^A�'1ܴ%� �u��ט�g}0�c,E�$OB�����c0�(x�;��x㍶��)�^�d�-x�9[�b���-ז�l*k�C�6y�6��:�;�H���N��jU��t�Ͷj�jǯ���`fwv~3ߓk�hB7����N���>�.��ki�X�z+�����'6�U�8x�A�ٱ��i礡�~;X�s���J�\B����4O{�����'_G�� [���S�WR�X�������U2��#�H��[���}x`�`�5��.?�/-PU,9� �@q,稜8�����Y[�8��(%\+Dk��*��{��f]J J���)��
urj��֨k�������Oi0�.Y�5���(Y����ܡ����h֠Jl]���U16�����7�D��+�(g�X� ���1���1c�Q
����lp`��Lj�+���w�e�}yW��:m��6u�t;���m�]����^f��q������En�F�?g��������S0C%�8��'���:�u6���z{�[kKp�6X6ko�_�Y_���P��~�;U�A�x*��BaC�,��niܿ�6�2/�H�M [��9�3�w�^�:Ná�V*��ŝ˪�󷦕FmE��7���}� �F�����UF'Bց�����u���@����7@3�:rfs�"~���q>���ǰ�P�$X}���.r�A.��i��qkP��AH{�ɰu�ţ����M\���o�;�� �[7RR�sr���Wj�FM�4X&��J�HI���t	�ׇ~�)�%@��B@��(��ߡ�O?�u64H�G�r-T~�vE��E��nc;ﴫ
���p�i�{��ahO�I[�H�k�WR�ab�>�;;���ɿ��.6}�v�h�y�v�i'������!U�g" 6�SO=�� ~O?O��)ڇ��?�����W�£X@d������
4I( 4:O|�V����<q��`ߏ��=+�s3�6���%�� ��ﰒ�S�$��|B �D�p/�s� 7���zA0�9��>` �1ψf	�@ @'r,4��s��\�Ǳ�[օ ]��m�X�xP2�څʀ�E&?	��9�j�2��ƥ��$�zR8w����	�>��B�}���������哀���� M���>hN!!,K�qf?3�8��8�o�� 3?*���>��{��z<(ԛ��z�ɧ���g;�8��|̳��|���}�1i�Sy��|�������Γpk�ʷ�C�'K18�B�謥� Tڴ�^g������Kd{xm�G����9�=�����#:�J�|1� <�lhLB6�/���������9�n��?�(ʹ*�K�s42�wM�R��ߥS��U`���%��a�3�̭Z�1�k����3� ���h�h�QQ�P�3����7�FP��$�?��5���M&J���V3��Ij��+!�)���q\g��c�<)����M��Ki��s�GO�I9�c9��4�kS�f��u��(��o��M4��$%�k��օ�O~��v�]w�~���+Y�{V����gM�A	P>�"�v�q{;��cm���9�-%�2tt��=��S^.~ͺ���*�vL	��dF7��gΚq���~S�q��s�t~�'��htͿ���R��b�r�!�'�=��͂$n�P�+�8������C(�����a���� �Kj7�=4�K.�������%{lb*�[aS�V�{�D�H&|�xw����"`�?��^�Xjr�h���������@փB|�+*��կU{L;q�k���N"����*�W�e���RX$|�'X<	�'�S��寪Y9��y�������0�k�W��^�`��0��2ou|-��F-�3�{l%�<f��|�U"�'^'�k2uk"~�v��; ��׾֕;4*��ЩJjd vS*>�
��P<4���|~�uw��|�$	��o�R[[(3aqo�Q�����C�XXmI|�����n�9fk�xQq��c�ɇ2@�3���dx>��N]s�5�9�}��j��7׊�!XDlLg@��������29�1�[m��ix��f�% d�|�S�rK�Yw�$?%�c��p��E}��qȋ�q�^��ω鎀�8�Ѓ!�������6�~|l
��>r�J��X��1��V��յ�@��f>��H�c�%��أ�:�kn!9�%P`В#�?���<QK�a��k�BeCoK�w�]F]\�}��KC�N���t������S�=����'���E�/�G�F��<jxѲs�׆j��˨�<��4�S �w欙WOH�������{.l���}#0LƆQ	A�	�b�VE|8Y�4�V$��=I��?�s/��v�2��Фah��Ѧ�
8��B;}���~����}�V�lGi����Р�0Nd�G[4��� x6At��8�3��˓���Q��J�s���$F��s��Xq�����߯��$�����f���b�������D��3vs.kF��a�0��^z|N�L�� �5Ф���y,(�^@>^�̔�4p�Ԭ�@Ŗ����)f��P�m���9�=��W���$5�j͉�1V@��/��-��ZK�
�|L��~�(���u�?�/��{Ml���%ߓSc�	>��l��R5�lD�Ol���i�M�?N36p~,���ȩ��� G�L{q����Eb
a���"�t4&(�[��-�������8xd�5Z�5z	E���B>c#�̜�<p�18�2!��)�'�G��<v��3L~��㇫e>��蚪���̋gB� (P�����<�� ��j��<E����B�9�lt*jJI�y��x&	]Yc���"�D=%eFV!�s�@"`�.���l�40��1|ox��Эk<�Ϲr�K�I�3ỏ,(~���o�A c��FBIyc��U�c|f��	���,�$�����w�ynRKsd���]M��9*-K� O�F��C{h�j�)Z��Y����{�:�+j���F}��^2�"P�[���E��O�<�|U"�K��><�B$�k��]V  �s���K��gNI(㧴a���9����"�T:��	8@�8��?I�=q�a"���z�B�)K��~�[���Nn��-�z%×h~P���Pn4�MDՉ�A`IS��r�+p��\�����O���Xh.CUP�:��Q*&�w5=���i7����+ƞ��	sc����x���6���k��fb�'0�"U��T��C�Ģ�糁y����)h]C�����1l�Z�i"h��67��Xm�,
QͿV#q��Y]�.�q/�+ A�:cD������.���g^T�pt�o6�cO/�7O�J�:J�����	o���d����Љ����Wq�����6�����B��f��y.��uyv :�s�.��_~i�Ϻ�'M�x�y��K�9�Mx�����j���P~g��x.��b�C�I�"��zI�F*ž��y����8]��>ße��Ev�-��s��4��p�&���ԯ����#+T4m}C�F����'�7���Fm��i�	���8�e����E68P�����j�-Pa�0@4%�H��8�
w��y�������/oX�Ζ�����$����d��Ҥ���pH����qrj��\[N]�<7��	ϕ0�W�) �f̵ J��$.Yrr��LkO݋��YJ�R�g	<���@�����}xO<;�������d�] �:Áy�A����ȓ�@�B�q.�o�w�8i�|/�Cd2š�Z�::s�G��"p��-�_*�C���}�(����3O�z\���W�%���4N
`.D5SNF 
5�^�~�
�1���wD��(�A����h�A&���K�!h�ld5��si�V��1��,l4=ř�@���V્΢��rP�D�/�7�m��N�F��ܺ�k��ъ����_��X����c��>�y�<�( �U�8D��&����̭曹��&�Gh�P9
��oU�Dx ᙹ'�����e��s:R*��15%+�u���R3���|b��L3�C��,7�A�<����^�7[�zUT	7D�[ �Q#Ifq�ŦM�nm�>��W��/��^*ݩ<��o��/�#���=}&z/����b!!�b�<c,0�	�f�~Bk�c��7�z]C)[� �5��Y��@�4|i��6��r�rY ǰ��81�R{��K� &��.�f�� ���t�fZ�,�!@	s>�	����|��4n�A�.m�EEc^x�>
I߇����?~�[J����o t�K������;2����X����,XB�S�>�g�����EY(�RJ �
�s�hA�N��O����`=���f���F�'` I�c>�`��#T�>=!�*�)8��Җ��l֬�m�?�Ψ����CJ0�D���t�8�'"�_B_�@���W�ޯ��	��[���sD���#��3g͸rb�z6)�6q��e-�ZN�@ҦT����X�\O{�簨��T�M���a6�;��@1�2'��M!}'͟��YX�i���኱�"EkH��Oir���U$��;]W�%�CTB�T�ȱ�N\�8%����Xm"}���T=�EK��E;4N\Ka|�uUs߿��Dhh��H�_Y�������xZ���3�|�s���y�=.��g ;B*	���yF5o��ǪDH�"+ �
���!�<3>�I���M��g��)�Ce�1��\b��GF,%O��޽��U��Ο}Ʋ�S4��a�n�������-_��È��?/�j*��p��֐�{	I	,�X�|m$ٕC���=*�r<�+�=���`�(	o��Em������v�Z@����`�y�v�I!:�J�k�V[Oo�ggs�����]� ����=Ĝ�&[�D�B� �-.���Х�iaJi��ڸ�X4A��:_Z����o�K�u=	�%=���_�a�kSmI�g\��3��c!!��g��������7��q����8t���ԙw��́"� w���#׵��3]	@�g�p��x�N��ܗ1�;�y\�.^�[�B3�;x>@��Pj���0� @�X��VD���
5��9�Ѓ�"o���5��D	8�6B�p������h���RY���5��/<��e8l�����<)r�'��%�N��qh��E�tl.�q���d<j�Ak��N���'�n,0�5�1K:�O��ϔ)!�pg`��AK;�������B�z�lhpО�;��1[�l�ku
��s&��?J��̣.���"b����\��h���c ��౳Y�4���-�A֎61 %kF1�S��H ļ��@�1�Z	��'�%�_�Z�w(������[C7�p|r�z��H 0l~QE\S@��XY<��=�9�q��:1�$�Psm>WY*�z    IDATG���{�
�^d������r�yzO�{��Eiq�rR���֐��|�;�i�|�V.�?��*[��n|����Y�~�lR�?~��n������~'���e݋��w�:s.g�[#IiW����X�d�c�M�����[���γ��	߇	��������������s;����_"G�4L-D��������4�a8��C��K�l)i�yY��i{q���/~�i��f�$�� 	��l^6*��hhp�t���'�$j��C�F��~i%��ka��9Oe$TZZT�֭�$�44rT�P��Q�]�s��X�m*�I�%�7��g���6�(�ሿ���2�f���ҸD�	����%�%,W�Y�þ��h ��<���`���@�7�Q�9�&s�0S�/�Pv|^�!���Hg:��k�tnSN;��3N���/a��J��(Mc�5nex�V!�Z���:��J�OL���)�-L�@N��E�*a�g�k�0�<� ��|��x�=QVX����9���;����K�ٝ��/W )c�أT��n���s;o�i��15&�EO���k�w���� �k�Hb^hlm�9+P�m���Z�}{��&d�����}�Cd��qt������I���
`�|�1�C(� uxӄ�Ȣ��8Wi��% `�'ϮD��;A�NDY+�4cA��&Y�L�"ekSIK��-�������L*8�Ѩ�bQ�A�4�ҋ���\BUVS���$ 4��?:���I�g�5M	%���<�E�i���!�_V�)O|���xM�9�N�_����GZqpȆ��e	�N}�j��p-�c�whiks�v�i~.�>p� g@��s�~���}$|e��j|�\%<�ȘB����y������,��T�M,L��BHպ��ح��ns�>�nO�k٪�7��:�t~�;�����ς����3N;�.����Q�`C�}�����?u3��6}�ǃ��Cl���I�C&�x	�㚢C(`�$#͗ʞPI4{x��_�E�ЬT$�x�����$-� �+��&���*G����Ǳ,T�?r�/�C�ݠ�dxg /��4�wBy):������f���{�]J���%i��1"��R
�$�%4e��/1� P�ঐI�ב��8�l�(M_օ�Be1�>��/IIF�3��
VF-���-?�,>�S����:V	d�{�Æ�/�u��3���.��?�iT��tu��=�(e��^Ƶ�oPl1奧YcJ�"�������z�2��;���D��ڿ�Jnd�xF��`~(��7_dS&wXGG��9���#�sK���
;�#m��l��P��>���ZWW�_��i2����3���|�Ս��X�l�]w�ٮ��Z�2u���d����<�+[�n��n���f���vԱ�ٌ�;��S���;�9~�T$��� �f�V �y������W�8�BZ��IҒ�*s\tE@�pB5�fA�*U�J2c��3�8�s��� @������Y���L[�c��Q�%pR2�l~� 'c��R�8�oi�G /�� ����ǪSct	'#�~��$��;q�S�=��+��se��)*��ay����D�`n%�@�DH3�Ж�Tm Y�(i��ro��i0���ޑ�QLX�N�̏��1�'��e%�]Y7D����;�_���w���e�"o�@�&��Y��).^�eoi�GQl��0��'ƛ�ZI�i)����m?s^=�Y��~���z����8�;�'�:�̳�^�T���h7��U_͒$'t�������{��6��-�gLJ����O�޽��=��\[�����`��q�-����U�l�̽���Z5	 �� ��(��g_�j�0�p�X �����E"ڠ�O(��Y��}Y4lp@P�,N4o>�"�cC
X ��h+���V	�(-�c�X��!�@)^�s���@ı,r��x>�%@����#��Cyj���A��{S�Ǽ6�(t# L?��H(�
!� 楱`��L���C��Q�r�ATcƘ2�*Ɔ�e�'�n�B���I�$�D�����q��K�zi�+	�f���X!��K�j���lHn+�J~����4��������ʅmʂc~�����Ip��!�G`̭, �7�Ǿ�={�����Z�E_�'�>�}A&Mj�� ���i��������v�gy�����q���zH�VͿ�̞3�������?�&ɤ�ɮ�Ϙ���������]w�e��l��EV(�ͧh�ۇU�cU[�v��=/��4��6��j�ڋ8r�E�_�$���~^r>k���=�� �?]����\� �hҮ�[� ���D�R!�A�@6 �6�|/��84��4{�� dXPb
��9;ƞ"� ^X�S[�����pGp�Mw�N^7��s�cm>�͙c�X ��+~zG�LƵDQ-�=��8�ZB�p��5�ye�r�1��!�$A]��;z�.���X��C�^� -
e��7�x��h��2#5b�t�Kb��\�ԓײ����y]�J�p]E�q���z��}]?��5�=뚦8L���/� ��Ų+�m����@����xɋVA�kZ�RM��E+��l��e���o����ו�{�C�6#�3ʺ�`���ȴ���OHh�]��?�{�*%�f*������t�1V.��E���\�i[���V�\g�b�.[gx�;rj������,�йP�3�I�������<�T�qj����7�KCf1�)�bt R� �~�3A4n�h@y@����;�	���U5ZK+���}i��>���3��{��#\�c�5[���ϳk�а��F�g\����b��������v���:4�l�XQ� �;Vt����M��jn��-?Ϡ"p��^ ��h�oE���s�K��N�g�o�%̽�L��M{�S+o �y_��~1t�
�y�.`d�# ���
�'%��[ ���Qx��|w,����σ:XÊ��3����}���`�ux��3ԟ�_��m�ݶ�i�;�g���"����\���y��*�zM���>��K.u*k��.o�l��Zص&����	M�t���\w>��F�?���g�W�{nx7K�.�g?���䓏�je�V�Zl�{�C͕T��u�ڲ�]68d�t���+��pL�����ᣄ���S� `Cv�a.���tg�Lhmti��4mD	iʘ� ��� 0c� ���f( �}�'��Nc��A��u�h��f)��}�B��0���1B0�q��b�Z�}b�I��-� ���(ʉ����k�D�W@�� ��;B� ߈�r�s)�|��=� c0�Z<'Y���.��� o���%�'�P�=��C���R�����o&b������{���w��?��2����p4�{��c�QV���>�яگ~����e�w� hտ�˿�� ��1��S��<�����;�C��Y�O�y����\���6�_�g�Y`����.��N�����������������hNa�U�o��Wv�y7{�{n�L�b^|�~�����c�R�׺V/����\��n]�-_F��6{a�:;�����x�ob6%�ڕYy�%�x/� �x�|h����O~�V��E�H!~ ���E�p=��j�9*��DE�<p��@y��@Bh�@(��P:�g@sAh���Z�|T����#@u�<��=��=TE��Z���O�TV�h8����|g��;D��S���`��F�W�NƇ�� Tm3QE�0WC>��������o�9繘/���،3�@x0�Xq�~�G�Y�ԍ����q/jN�Ys��P��=h��p4��p�ui��ǅ�t̖Y7�s��Ϙ����v�[|%���͚&G��o�����H��8����+���ڡ�c3fN�^���2�A2W�����-�r�Ŗ/�[�P��|쟼�iw�:���sYT�4��̪��c��/t���4�Jp2�������h��>km�ط�u�w�V.���e,�_k�����Z�Ζ.]iUk��K{m���eeX��,�h���7|SJ�C{@+���˜&��i�h�z���XXrk�� /�f� ^�L�C!�h���"U��o	�)�����������[|��Y[��u#�5��ⵡ"���~���M,���c��������\Cxa�J���-��y@H�G9n���x��k��V��Q���S�;j�uy�)kQ�g�y�x��!�'�h8͕H)&��-���	��	������ܷQ��%�K�"?��k���~�aW�k��C�A����(���J�͟�_��9{����C���۴�s���P��R��E֞|b�����_���d{׻�<��*��>�9[�d��q	>���c���ZҤI��w]o;n����`?���e��T���k=�~��,؋/,��]�mmw��?�-^	&$��~%K}�c��s�=�Ԣ��E�H��;��/[��ə�8�F_�`��I���|��L ���EI�i��t9ͅk�q	�Pf�d���Ikk-bHQ@�6����; �u��I�S<~[Z��{���=�??�S�9+UVL|��P����!h%��c(���z�}���a1��b���Z�2����\>S�#Ń��`�<��(0h���j�!�>t���H'	������׃�蟗r�M���;͹|=��1�>ڵ|.�h$���ކ��j I¥�3��V*�����ȦOk3��k�J�z�j �,�j�y�X_�Vuu��g̶SO=��i
eOo�֓���������[�\?^�tG~)C��?�Y�/�]�ٙg�n��>�z{�Zo�:[�f��^�Ԋ��X�
�P�����ޛ��]����Yg&$$B"�B�w"�Z��IP����ź�o�׶�����V\��KMX���(UPA@�%����6g2�Y��{?��̓Üs&���f�����[�����7R��n��$���]^���Z��c�5�h��[5�Ź�lX�9G�K(��}�r6i�*�`S�v�J<��^��xnv�h�C��܏�b�'�h��{	E#I��<�T��V��'����u	%�8�ǻ�X�����L� 
�8������	�J��w	͋�8H���w��%�]�KBw北�:�����d%j�c'&�AQ;ʚ�w�}4ǔ�@��Dsƻy"�~Z��0���N���(��yz���������/E-V�� ���Z��S�#ʕ��E֘�%]P	,ٺ�)۸i��ض�JղM��[-�����lp�j+�Zk[���eo}�͞}�U��~�;����l�#s�h�,��_���
��w4�} 6p�Cgۻ��v;䐩V���y���l��uT7������������C��N{�2����>�X�;�0��+�ʿ�Z��7����/���f��6��s�Øwf#+kT$�H��"�A��7����'ϣ�mi�Z�z�84��^�v���6)!$s_����eE+�~��������VA���&ca0�H��#�� ��3h���w���u�ݩԂ�c�'��X�`.8^�ɵu��+s�υ�������<��k=h����]�G�:��?~�;��W ��E3����������G��k\Q�����̄�rX6@�Y�YG�j+W-��+�yC�O2)UISV���u�y��c����`9���o�b�Q���V#�Ϝ>��ŋ_�8G��5�|��Px[3��dj1�ɋ^h/y�mBg���)[�z���w���k���-�-��ڬٳ�����{�M�p���¡B�P�MY}6�e����͆)Φ*��/�C�A�C+��6��ٷN�H�i%[`  ��x�7�V��.��K��I˽����J�����o��d���w���v�W�X�I8�z
���9�o��OE�$�~�Lڲ� e������" �oqss@�#�j�K�wZZ�Z?z�V��-�+Y\�x�Ю��s��Oi���9�_,9^����Z��U�,z�}4�d$���9w�(Ǘʡ�&3��L:G]����Ю&�p+�?������}Bg��c�s#��[��=��mdN����E]d^�r�V�^����,�e˖z1��g�9�y����̎:�y�7���w����Р�}=�}���;7_w�������P���f�/P�=U~�$���KmE���P�3��߱���cƌ�>�^�;���l����YX�~��}CSo?�'�E����rE��B=y>ORK���QYh�W���?���;�/?@��wh�X�y�X��CDE�rs��CWI��i��(��	�h�����|_�?�'n�g��Ϙ��V�Vi쌯Jr<mc%����s��BSS�Ɖ{ro���+��9
�9��^s�8�.�*	X渝e"�wAc幜���I�B�B*��y��Z	�X IK�����Z�\��|βD�O,������pP�J-��0�����)۷\Jh�&�ߘD��.<�T��h<��ݗ_� ؃zn�(� �v�*�%�O�l��vt۔��G`��#��b`����Z5�wt�����?�����B���'��?0�����.���)��w�PŇ�r����7�ѝb+4�����+&tǎmo��lHi�L:M+�� 
 ��[��V�U�`3�~������4�j���b�1�<<?��;�#ԏ���R���� Y���Ȋ xV��h�h� ���(�#\ �����w��g�TbB��8+�������e#K�f���bR�f=��k��}��)u\�1㠕ƈ�!��3��zH*zǆg-	LCƖ�b.9��C(sՐ��J��J� Z�"Ɓ
�D;�7��:4s��o~SO|��P���t�Ӻb�.������{�΂mZ��K��ё��M�b|�?�Z(��1ɦΘi���\���~���m��-�t�I�3����+h��+%G!��Zan�3{�t��"����c��;|/֟<�Q>x���e��X6�	�lGֺ:����R(��u&o�����?��;�Q<;:r������>c��nY��+��ߦ�c�[� kq�c�R����?����d�׿*&�����ʖ,y�^�%v��G|�]w��ݐؼ��ԅ��
��G�v�-A&�q��N���zQ�@�I ��ffa�0
��w�$#�k��.@Ģ&I�Qug ! _�HBR�H��
�8��1�t��3�q��V4Ҿ�}ėJ����:V�q�Xm���i�����T�&����g�4�'Y��	�)T�XT�[IZd�2~܏yc���/��a^G�S�Z;�Gt� n�e/{Y�i$��G�+k��^��C����%!�(%��sϱri��{�~�*���\&� �
��ZMp=��'b��Cմ�>�X�5k���6l�b_��{l�A覰,����#�u�%M���.�>s'kPY��Ε��P�s���<���ʎ:�9^I�=�N�c)�LV���ݕ�L6������ZP?��߮�;#m�IS�~�-�|���>@cp���*Ւ�\+S|q���I���|�	�I� 2|���x�� ��-FE ({Pe��w���� x��&͓{ΊL@!	Iڦ�F5o��`I ڪ������Pb�Ҍ��І%(��c�S<����Yisc��|��u��[���-򪬲H�)�ڌ��=O5c�Y+l|��f�'ƛ����an��5�B�C �@�ɪD�o���܊���=@���*�����P������������[b�u��V�Zi�6oXo}=֑!>�b�r�i4M;r����J[-3ѦϚm��j�j�
�}��k��ǟx�)��4���E	�� ֘񮪃$�]>1/���7�@F@��ɜ����#�������p-p�`��g�Ppq�[\�#O��m�f�*W��w�C�W(��UK���������B���>���F��
�;�x�5��    IDAT�B�g5YV_�R�/���2�/�i(����O�����^;Nk @$������rN㚊��Bi��(0�f/�Ţ�z"��De�*_E�x+��H�q�𾀓|	��POT�~W�6ׁ���2�5`�;C���{_���~�O�u%�>��@	2_rFs,Z�֔@a$��Ɗ��'|�o*�J��7��]&�c����r�s����]-�s��'�Q�xY	����?���=�[�@�M�r���w����趘���Q� �TyЬ<d�V���7[�Be��[��'/��CCUO�*��Us��9G۔��:�wz�_�p�=�d���!l2��.��b�Xrq`�LD�%�}�}�K_r˝r�u�]�E�"u�1��͘8U4y���o���PV^�*�?)��P�A�w�'���#��6�g���)�����=>��t�~ܙ��ģ+ X,�P��j�] ��OX��~��C��Omj 0a�Ӳ��f&���}��"o��3�i�5�U��X%�(�H}b�q�Qy5�V	e���`��,P����Uw82.� ϳbEȼ�;@�s�O}h?5$G� �|��/�k�\�Uc)*l_9|���i�K��&驿��#��
��8w4:�� p��\��^�U~�VI`Mh#�S���3�|�u&ڌ�#a�Ԏ�Q�'ϫPN �P2@|�ִ4����J�h�D��+���s���{,���Ƶ���c�ufҞ�J���~���8 תVM�l03��3�&M>���i�6��_���VZ'J]RZ=r�֚���|<ק?�i{��<�| ;�r.�k��}�<� d�3�Y
R�<d�X��4�D�|N�"~��}),�5�ã|�7B����Y	h���}*�g̼�L�j	��M��W/_$9,���31 VtO�P ���*�aP����������y�Q�i7oݭ�U��I!ڠ]��$L%TR �������� ����DkDp����y>��B&�@����;4Gq�,`��g��:��Q)��V�R܋��Se��K�_���g�]c��͏S#�q
%LT*�;|(�h�|���YT[�8�����P�*��5���fYc�J�MF�h�N\i���M��%��=�X��
�][%z�K�0N�Ԁm��rV�5�V��-����Ւ�,� ����TΪ�iv��ϵ��DK島e�v��k׻�c4�����?�'i1�j���O~�֬Zm���7����~ʂSߟ��1�Þ}}�k��D]ʊE�ↆBX1��I2����#���Jz�|�O�V�̘9��o���_k<�}����,*t.Q�'��	��K8�Ɨ�$c^�b�[ȥ�l�i��f��|i�, �8\����1�i���f�������s��sU�+�CX��N���1����E�v. �'@��@·
R�H��X�*7�3 ,q���� � (Y ��u�w���x
��DК��G ǽEY�V�C�Z�[\9U?U��Z(���������{	��h-1?qKF��|2��sJpKH�* �IDOi}J�ig9�{Qh��yN���i'�`��+C�~��c^�����ͤ�����A���?q�A���i�7m�k���=��S�'YJ�kY	�4Z͟{K@�;DΡ�S���N�(��0'�7��/��/�-Z�w�Y�A�Y򱐕BJ�N��)�(7R�5�T
ڧ���ߊ���-�I��a�g@��ed��ؑ�zh�f�6rp'�����l
�pπ�J5��]K�KE�p��.�f1�%\����z��,�&��k�+-��%
�N�)�x�[	1Q^zY>\[��! >��w�j�tہ��~��k��ߧ6.�)G�@V`�؈;����A|/ �z�
�JK���{�ΕI!�����R�RxX#G=S]�%]��.�x}����x.5�܃:Bg�q�k��r�i������W�N��.Tm�6�τ����߶�`_������K�ӹ �{��+�_�_
��]�� �1g�ׯH;|Z̟�nY�Z�4��A��9m���8vi���@5,�)Cs�j�[p�8O ��	bT �2����F@j�6��9)��'<���:�Mh	���L;�ԤM	|���:|/� ˃��9��:Ց��Ε�(^�Rڹ�M��Oi���j {����3~�����������v�Y����x��4F��"S~[e
�X��Kc+kP�1fXr
�%̹����@V�"��%4W$F����<�-��;�z� %��8�T�Ҁ��l��ֻs�u��CA=�\����;X��G?�&O9�JՊ;|���km��-MYD����h�I�/TJ{Y�1Zl5s��B�+|r��}:L�p�D��ĉ��aǡ�M`(��aއԑ��8���n�&�H�x�w��'�$uК[���~
��EݼM4yi�,8w6���ht6�6��G��1�h�I𝀸t]I,��2��'�]i�a�,:������������g�<���qכ���5��[�RG��(�4 |���d��=�y���%KB�p�rbK�yD`-p ŵ]�I��@?^��;vr{�H��²���Gkݶy�-�ԚC����gX�<d��۰v����p���X�])��C=�ռ~��6��Éذ-�wؿ��ڒ'���	�] ğ�̓�	u�g��-8hC�����+�H{/�S���Byaܓ(�B:���q*������<��7[��}�å��,�$��'��A�%����Z$o0�[�n�|E���<S�x,xb ��'��Sa�X[�5���y��Z��b�ǀ��γ
D���Lև�_����k�1xb�ƛA�I ��0�y&(�_�>�<�1��V�A�q���X�J+�/f5�r
�u� S�R $���� ֕����K1�wAP�+���V������4�����M|�YgZqh����n�`�};]3�=��}�zy�9N��6���6}�LO��oL:\�f�lϱd�j���)�Z�{SV����֘�Ա%1]Sub`!���+K�-�,�$A��l�q�g�U9a�8�����3�N9�6s��I-Z�9ߛ$X���]i��9�L��� TG(:=�|/�1��c��5�H��4�F��X�-Pӂ�~Ah��&-�V`�0��5��Jck|T\_QJ������#M<�}bMZ=~e�s�6z��^��K�Z!v;�hT$�֐Rc��<�^��敟��@9��)jH�C|s���ח/G�+%{:��x���8�=�7e��;�s�\����?�{$��p~���/�L;�&M����t&�͈z�	�{y�x]�oQd�?�B!�!<�)T�$V�4�u�<���%�v2I�"ǖ� �#k���Z�|vu�����g�w���74����h�6�_s3j��OU��i�!Ty��uV��qG��	-�����v�g?,��Q �w�7���s��cmN�/KC�F ��,J 8�2����%bm/�$F2y�1�Ij��D;�D���p��]}-#Y-<���B����I���S��4�=�UP�B0�!k[m	�T�:귣���+��w ��� �t,e/���;�Xo�7$r��wYd�����w�q�\�g�6�Xu�O�g��?����Li7V#}����֑�oϚ/-�U=т��"�R����rŲ��l��e;�Dh��YB��aa7)B̑�]މ1�
e�Uԑs�N�_�ּ�0��lG�[n$l�P��;r!����CuR���X.��a��V~��X�o]�!h�>95����7&o޼s��Shf�8�7*�*��v����,&Q�>ͦ�?����c���wo�Q/�&-J=�x��ħs��?QA�P�֢��(��ck MK�]G�[�}�����^���zҤ�;O�2�}M���K�$�s��]*$��*5�ԛ���n��;���@����_Q�� B���o�ݣ|h������������A�A��AV)돜2K�l~��_y�!�{��_�E�PD��d%��q�����T����	��Z�W��Z�����%�fRV���9��V�f%�}���Ý�MI�0GP�t�J���aI瘮��m��J��+E,Vd�/�r(Um�DҜs�Qv�s����&L���*p�|�
[�jm��9���wtUUh�ߦ�[:������zgʪ��o���E6��s|B���r专�R�y�Q������M�;�(F�W6�w�i_|��� n��f/�,���B���&Y
�}L�H;�ƌ���v�V��"���.��G��o�L�*$H%��]�P7)������J���4�%#� Bat�g"ڧ�;P�3�$��'���_���l"Q���44�v ��ݾ��o{���.��rX�4���_^_G�]w���34a\��^�'����?�����ČG����g����̥qݱ��B���̕j=i����[BC~�u͘q�W��;�8�y�t�|����{����k��ҥ���w��a����;���g��i�r�j�Z�>c�{oY����u����-4������P�L>lj�ܜԩ�_-��n�L�^��/8ߦL�T�����n%�~�͆d-Kel��^��^���1@S�����\k#&�l?��O�/x�oR����ы�Q�)iӇv�&;�H&c�s������Lp��( P.1>�`�w��OL�	���X3���{�񓟺P�v)�E�.�&1�M{!5���a*���E�A} (����J���??h�q�>�nD%��CH�������3n��F�S�r l`U��J(X	���Z�b$���7�#X�?J�����|��|�7����b]q��y���BG�&�\l5ǁ���������e>��H�ճ�/^�:[��'ͣ�"X�V,��Cfx��'�Xj�/�D�\G�	�'	�#����V��Y|�^B6oC��v޼��k_{�M��e�tնm�l+V,�%�?b��l�,����c'�x�}�s���ȍ�SA������/4 �۩�����}����Q��+��K�,�ו���
HY,&z�"@�8P'�W�d%����v�F�l^�W� �>��j�/0�3���[ns�U��w,�Z@���)��wн���)�����[֯��3|G#X��<�ǀ?7E�����}>��	�#�i�A) ���0(�} o�h�����6�( (%� ��J,�������}3YN#�5�w���Oh�.���_�}�dK9����U=|QT�O�-t>���4����VX/eֻ�y��m[69��!3���͵l.o��Xg�{j�*/'�z��?�h���j.��_��?
=�����3h,@*xN��f����J�1}�UJ}�}�f{����򧞰����iV�x��!���?��<{� 6����
C��_�����|�+�G#$=�]W\�<-ş����E��i�b�̵`�7�E�l�V�C�����_��o%)�`���i��Q�	�"�~l�[n���q�u�G���FZjD�#m�����?vFslɆX����G��\�5�wu.c�Ӵ@F ��W�(� ������d^o��G�G�W�.���_K�g���w�!����*Ҁ?��I�0N����D���O+��{���"�u��g�������÷���>�N�G9 ��Cq���g��H^c=#�����g}#�K�?�7�\�Ry�{�a��{�9�Dp��6�?ds�e�}�͞��x�G1��n��P
����9���M�r�8��T_�k���۲��-y�!{��-��zQ|fY�e�lgϠ���q'�j��z8ߗ��e�p��{�s����I�OU@z���	ƥ�H״-�F����"t ��5�q 	��f�NL-5�rů��*���B�i� ɢ�;��{�}�����K.�gD�yN��IS�ZV�,�}�9`�{�+���gV�Z�w~��c���9����p��O'1�D��{����h����5�s��� a��������s�T��5��;�cF��so9|��C���D(?�e8yk�>��p)#�1�ozӛ\������[xXq`��z%k���\���sө�elȖ.{̖=������i塢w��첁����؉'�f��y�z�,�,��f_3���4�����k�N�6Bg>o���]��c��T�h����6uY{�l��^��R�����l��-60h�ik�����y�?&�g?��kq��1� L�/~��&4ϸ�7���dS+$NL� ��9�|�T����88���� ��^롃q$�H�B�����1@?|4e�#�U�(���h	!m��8��m���?��'��GGçp��>����zVǩ���G5�YNz�/s����8��P GB�n lE}iޕ��#Q5�&c�H2��(tX�c��q�OE�R#�۽d��u�gl'5��u��CNH ~rB-L�o��?����������h*X�>�j��p�c@����f������8�k+�z��%��ښU+Bu�rj>7�֮�d�}CV���-o}�<m�<���d?���u!+ 큫����U\�3�����:<�䆯~���O�\�+��_dCfҝ6�_�IJن�v��'{�*@ʅ	_�0A6����*@,�0A�C[ToV6&�P�D���׼�����PWg�h��.\���V[�xbU��u�<1M�E��_�!��K������V���p�bR�$9���x'�h�h���sEg���
e�. �xʿ��}���.��r�_EH�Sf�d�i����u���h����^q�hȝ�P4}r}��a�vCͲu� ��m�\��5s��w|0�l�ga�`�C��/ Jڗ��%�A�p~����ۻ�CgL�I�'چuk�FQ�u��r�f+W��J5c��vۙg�k�{����k�-]��n���m�������T�s��q��?�c��Q�~۸a����;l޼S,�.���Ox�_b�k����m��V�u����l�	��#���&���|����	11�x �-�_����:�JQ�Y� �Z���(K0Q4\0@����<M�@��qBSi`������Y�ȝ�q���]}/��������D�ƅ�u��1�{�IJ������<��T�����d�ǚ�(A���c?.���j�����Bz1�-KNV�֔�Y���؃�����E����$vՂ �4�g�c���aܘ+�p� ��ĺO|���u��,p��"�/���l�#��_��N9�h�1�[�أ60��� |��@��u�u{�uvM�_�q�wM�����ƛlŊUu�����p��3�������o���>Գ�毥v�s�t �Z�V�z�~������n�T�֭_i�}=I�D��-ڪ�i�m�/�`'�r���M6�wh�C>�4z�^ >��?�&'�mTB�LR0L��E�z���d����q8����Z��Z����+�tx>�Ef2���P�lFۇ�G�W)�v`?ҳ ��>�J5ǆ��y���P|�`��)���� 4�틠m)�E�)	7Y��W��9�k�B��6�Iܞ����z�XP�^��i�~��n��KV��^�*[�x��k�c_@���o�i�J��;o���8�>x��Z�<�zz�0 e�=���Ga�v�����~β�N����o�b�r�	Qy}Y����?_ڬCg�'?�1+�,m%��o�h���ݶy�:��� S-c=�A[�j���Y۸��iej��ѫ�O�����L� q��lp���7;��������ϙ��)�ub�w��A|���3�n�k9RZb+��H�w,_zH1�#l�/>#�p|�a��d
)������s�|�|4�ǳ���c�Ɖ^��k�ɇ}�u@���k�|��������5����N��`lEi�]�u�N��'�G��6y�Tۺ�ە�U+V���	l��������w����1k������i�{���}�v�
+��i�N�mg^��v��m��m��ګ_�jN4    IDAT�z��=����N����F��w^�.����)ޜ�"
ɹ���8��e[���L��4g�� J:�xB�	x���?BVj>��Ku�#�>�x�!�G�/*N91����N���������=�C�8�g�b�;��{�#f�Y�kV�p �8���oK�\a����M������ezh���k��j�=����G��V��τN;h��v��U�Cֳc�mߺ��wo�Ri����%ˤ��/tÆͶb�FK�&�;�����~��1�h�$[a
����O,�,e������׻U��H��J�#�x\��}�
b���8rM� I��~��	��磈'ێ�!
��V|SK��n�������ڱ�{L����C�N��X���O�Mq�*CQX(~�;{�R����l˦��ݽ������}#,c]�{G�=��%ֳ��.���6k�l�T�v�O~j?��-����)��%cx�:|���QU�t-ms�εw�������[��=��a+�l�L�f���@����c�©6�9�8@������$ƟJ���DD�"5֮_��f��0��deӡ��H����?�m=~�31�p��V�+ �Xxj�  T(Q�s׭�����G�3!���c�1�X��V�]��ʏ}���O}ʁ���\'J��N�qQ���8�@	�_�q�h�V-�e˞t-ʇ��\�_���`�N:�t�{�)��uX���]��=� \j% �8�VU=�VO6D�,���)S�S����V��k�����k˗=�WS�5a��z�iv�9���鳼�@Ov%�J���D�/Z	�-���� ��N�V����J-s���7�5d�9�q��X�l�+�EV �1�OTq(t��1M�HłA����9���,h��<�x �XޓwW4�"|ؓ���<��x�c#G0>u{� }@��˟gR4?��=^t��T��Ѐ=��v����+�[�J^HH�<a��v�ة���5���<��gw�ү����s`W�lQ�_]��JE��5�bG�������Yg�n�Ҡ�je*؎�[��[��'|�t�T�e;�X���y�ų�0�lU�'��/�ω'���]D�ȩ�yh0,.�>o�1���h�fe�h���]���3kmK����=���TB��b�e��T�#�u���Z!����eK��iU��ݳ����Z�]�I8�	�&��g�P��������,E��	=����ՙ��ނu��ڵ���c��>X3gf�"��t�._f����~ *��Ƚ�g��o��Uw���(�J}��|_����/8ߛ,PB�hRJ�ԩVC��޾�����=U�/����W_�@�ǂ���+}�X����_yHQ
,���ĉ.��9�� �������0�S�-�]�z�gvS���P�b�W�H��0�U-�N۱�k�$B�<���z��р|�cT�	P�ު�p����+��Q��`�<��Hй��P�^������_w�[t,+��~����o�B��G}ܾ���Y���^5�\�~?�����
݅KGN�ҿ1��o�P+�F�&L�I}��W;mCyg>��eaB�l޼ս�j������1hj�v���A$;�ݮ����¦�|���f�����u��E/��pdƺ)Z� r�YH�m���RI�K~��a3C�ocl��Iy�V4��s�єw`̈��Z�ot�kG��hL�	5T�ߎ���l�ќo*9��7~/@�3�UnC�[��O�c��*˺1���F�&�4@�������Y:������<P"�s��@V*�uMԏ*�����^U�U����Ο��:"��G��t\��ڱ`b/S��w��l ��_Ia��vK�N^ټ���!�ε��&{73U�,�"���3"���==Ng��O�������3�?�{U�er�w ��9�|SQv�֊ ��kA�����z�^p�c��G�'�hB=�N \i��$���MD��JU�z�J�1h?�z���ΧV�C���0S%yQ�ᐩ�F��5K�P��| ��H���I-s6�j��o�AJ9��y�X9�v���PVl�Vr�	���v�h�}�{�kK�� 9�5*�9(*I���<�ϕ �2ʄf?�0�}�o��"⪣�KZ�?� ��GQ�\����C�k:�=y�s	�x���8Fu���
#�{���zdN��\=�����I'�uE��1.���}^��н3��gýR�`!��F�w;����߬\����!�������`;�Yw8�� R�l*d䖂êqQ�����'���� e`)���O~�K1P��k0���Ь�Z����uY������/��K<;��z���$�8r��w�'�2��1�uI��nu�������f;��X*!R��#�*!�ZD��9����ƒ{��۝��R�S_'I��:�\IJøގk�{��%PdQ�Y���M}�����E7V�˳���R*����7�(��8�X���r�����%y�w�q��ؒ�] ��v��|�a�8�9����&�KR���_ʹ`���Ă�n��(���;��2�j(՜��10��hh�����©q�aځ%1��W:�����& ,��iQG�k�$��(
M��.����n�4��q-� ����S�3Lnh�^L� %�<cA�CM��%%,Ne3rV	��B*Z�#-���H���i�����4��y󭷸�[%k%�)M��c���;���Jƀ��&�*�;�I<��6�~�r�&�����+n��F��I��=�w�y� �`Zq���)�����gkw�-��땠Z�$9�S���Ny �͟�J��/>88�'�h�=�H߫���Uq,悬b�Q��P'~R������:��4*�uKh'-i�T�d/�I���z�p��`�9t���c����[�a����:|��)�<�n�jA�G�
�t��b4�J�ĭ�r�w&NG/��D�o��w�Q�4p�	��4B)8~B�`�?=}��\RW��O���P�v��1�ƢVm�F�_�E
��@ʂ�7l,0�	��ӤƋ�Ն�����8|���t�Q?5~D[�n���$� -���/�_�\��o�y�V�֧�㿧�6�S\��)�d,��1��3>�C��D���1�ז����+�Hc0�wP䞔Q<�p#t>�񏏘������j�!���ZA$��t�M'�%����.��{/&��?��S4vj��9�ƨ~��0��̹j%r �p��TI���F팉Ŝ��o,s���v�]�a3�q��D#�����y�E���c�G�̹^��_���GE� mC�&	o��%���9|o��mN��;�GμUO�}|���ռ�, 61�<
�y�ERu�&}�1	�?Pn�~ 5�6�Nh !�^c���7���X0�bJ�k��%81VXI��sٝ���c��Z��<vXJ��6�ؖ���5��s-���}ޑ�Wt��>��{����M=���s	����#���[*%��L><Y�h�`����j�P�8(��c�lοE��k����HӚ��L#�j��PfA� �Cㅴεهs�h8��f���3�T�.�A6h�Ī��x�K_��_o��ݛ|���}ڙ�.���K(�H��_�����YG��ӈ7'�}�[�����Z�%�j����p��&��r��`����(��7�_�`ų���ʺֆ\H��Y��]Ig�� σ��:�hr�]�!a˽dep�7��u�[k�v�DϠL�՜�=���/���Z�7���/ņ[�ַ�o�(�MhY�g\v��۽����u|/�E ��Ou���]4
3)ij(q����^�B8y��� �]���B�'��F�g}�}�$�V��6(��������J9h"����kv.�E�*b3O� � Z���j*���U��lp	��h���z�����k�'�3s}@�{�N��h
�-	gv�Ӝ��J�½�������v��L�,��rSI��	-z�	��d�k�	,�m�=�>����
��y�K-�f��ˢE�p����ޚcͫ�|���3��:�_|�cu
E���<�p}���{�ܘ�z�K]KN/�����|
l5�;�m�Gćs��#k(���k� 5�w���5ͳ�}�� �@D�����}���,��U��4r����a�N�c�}��Ĺl	�f���]g�aV��%���ש� Z�j�qԹ,�봇4�X��$���ڔ�`k3K[��N	��G�^���":���7��ɤsP;�m�X̭>��X>ZԊr�i�+C�N��X�m�ϭ1ֳ�����Ƈ�cݐ�G�a�k���W�q>
oe^Y7$���_ �O�'��ց�ќ���F{���H�VS:᮫� �(d�1�K���G���{�ð��OJ�H�5d�"n߮��j�����5(�_ᥚ{Y$z.�����)+V�\:��[�:��0aP�p��q�R���bZi����Z�UfN���ŋ��5�I��z\��n8\(�Z�f3!<m?PA�
�d�<p1o�9d�2�����[2��P|���^��/ ���r���AlA��'`�l�*D��e��iNc`޳��c�T>��9d:k|��~��e����{�U�k:�~K�.��2������C���x:LUX��|��zA�v�/���g�9����E��e#ϥ������+�|߯��u�^X�-���W8�j!J��s�,)*��%�yX#t��3d�Ha�<�Zk�fَP�'��Tj�vM?X��/���l` 亠t��������fQ'�_�iH��gsA{��ET*A���	�삏/�dtuM���m�G�X��Y��5�"r$)����`���18�`k�O����o�������c˪����6
���v�?��ey0/ZC�B(���ؕ@˩����X��<�@D��Ɖ碥���|����xʊ�T8��=��كs�!��}+�_o-�.�ZPb�v�':_�[��["�CG������mw���g�a�C�JV�r�k�o�	C·"ɔ�r�c���OP:�Y�Dw��f�h,;�����eѢ�5��[��2�vH�pS*���<ҙH��#����zz��9��*k��2��7W�?G����i�P���c#$X���A9�c�kԲ��Z��z��3vJL_qSi����3n� V�\4�.n�'�I{$��a��r���D	<	t�ݓ�.}�.�5XG_�����+ϱ>{੓���[N�Ш=|����,���-T I�5�kX�D�L	����eB*�sR��E+A�č�[�#�	в���i5t�#�PX~ �O�?�"��-ʸ��Q
�|H|?�2�}*�O�4�'�@`��P�	��3�-4��#�wIݓ�u���{����I�ä��j����+��+_��L�4w8IY�h�ī��� E P�����P�Z�5H����t�Ӥ{���6w;�2Vڧ�{����힯����^f�45�9"����ii)7ɉx��7�R`�M��m6o�E�p} �� W��}^J�gQ�I4j�l�r���+�%A�t��(����^���{��QC�lҫ@'as׸��e�r{�q�^lq��aD�o��*�u��-<�,�o�%�޵�M�4��e�E�S�vJ���B�ּ�1��=���g̜����{�N^0<�=�Č�8a�k�z��k�>}�o.����pg"���r�
���d3�������S$'}�{�sm�c�S)��G13�Ac�yGF�D��]�����H�c�v�>���>#	����{����Ώ��;�M���T�t~�����Tkgo�"�ⵡȣ|�^AR�	?Q(�$�Y���a,c[n�3��ц+f�|�.�G�A��E����vy8���o�����w� ��h5�/zE��
��=Ĺ�o�g��	����,a���7��N�����3��a0��7�a}�\,��_����w�s�K֟�w����s`g�.���B��f�?���W��Ͽ���/�x|_�I�>�>��p#�-]�G}ԋ�!��X��$/!����!d�&�DkPן��4|�\���`m�FN�QP�u����p�÷Q���tO�c�v�����������d�b�1�lf=�z�{��^=�}��6����@��8�����J���k�j?Q���U��N�8-����9RO��:���^��:�SW(v�c�˾dL��ȇ�ͬX���	����n���d_��?��{�'��"�:�'|ods6y�A�y�6�ݸy�w�A��r��B#���m���5c�R��l޼y6�E^�&��o�f�
Ϛ���O:�4;��6g���2����#���7��<>���C���?����?���Ԑ4 ����E�&QO K��'5�ݱƺ�������C�'-p_ܿ�5�PX+hb�����x�����$�v�s4��2�&`"��}�)?��=V�����}/�Cs�s2Vʒvn��|
�#<�2�I(u��'��4y�Y?��T�z[�:�X�`1P�ΡW�%랂����~�m�C��W�%σ0�3��/���z��1����_�Z;���B����mt��rQ�4�����$�;\��Kig��8��3���[�F�$��Ϝ9�.y��v�)'Y�4h=;�ۃ������>!D��P�{�̙��9�γO<�r���o��v�Oux�I%J���ϸ��`��ٞHu�M7�BQ8� B`o�v��@��g�T�)vp>s���TH�Q����k��ۃ*2{�;�a'�=ޣ[{{lӆ5V跮���xJ�V���� �P7%���s���I���ȭ�
�쩕��uBI �	��s+�K|=���uS�����\P����~����Q�KKz(����g�A4��fO<�����_ن���EG�;����K_�J;�i�����3�����X�Ԟ|Mn5%�I�����=2gh�^���eo~����X�V����Gy �Х,mIĠÎ�ݶs�l�}�)�����d|�_p+�L�^ij�	��B@K 9�@	"\G�9ƪ9�������h����}������ڶ?%�N��J�^�nmw��|���:f|x^�8�qکf����{mӺ56�W0��)�x�\y��@瓊VLuج������X:�a�6o��v�=��ɤRR'��w�e�)���UI/|+�X�m�v����*��d[�s���N���?�K��m��'l��mǎm�ˇ���ض�������/p�'yq����5o ;�������G����f�?!��\Ʈ��]v�	�[�<d��M��a=�M�a#NU���P�6o�j�r�zz����y�{��o��>�
�BCIJ�FS�o���1�X�,�}�����4�i\��7C=�=�Cy��}"��Ya9��Z����[��P�m^�����[6U�t��QT~<�<4)��>ڮ��N�YGk��l�|�mܴվr�W폏>�+�N8ޅ�nr�%j���|�9�9���|��������+}��"��p��|�	�ʨ8�g}=�m���l˖��}�V+���O~�P�f����[�k��v���d�Ϛ�>GJ�C5������1��/�����U���#f٧?�I+ؤ�v����K_�+�ؚ�O�P1�Ϥ����o�W���!�������h�+W�ts�E�v�$oȞ�/QB����x!��(7I�g� P̡j(5���������)��=j
:P$k�}�{��u��V+Z�<`�6���m�,[��UܑN�r�g5�\��8�	�TƊ�)v�Q�ڄ�S,��t���7ڣ�?|4%v�ǘ��2�����g�����'?���wB�����>g���o��(~D"  �t�l���;��C��	9[�f�����~����mɓ+��s�-}r���%�_��I�z��-[���4�.92��`Ⴏw
ok�1�s�e������%۶}������i�t�֮{���{��e�����    IDAT�b�o�������csO8���	��/���o�' Iߑ��kV{$�LH�\�7�����G��J�ߛw���G@�}��Lo�P}6Γ�3��Ph�r;��ӬZ�L�d[֯���sT���x!!���:���9G[��If�[�q�]�MN��5�p��c3�PO%g�X[�k��N�o��o��ˇc��K5�T"�pN�İ[���_���v�I���i�l��%68je��R���\j��D�)XG���G>�e�=�._���ڨh$��f̜��3���7�oo��cY�l�a��UW}�2���Y��������ϰt�h+V>i��`����m���f�&K�'ز�[�O�+�����p�0���D�Ш�Xl��p-8@��r ���`e	s��8���z����N�V�K�z����1���Ͼ`ݣ��š�rѶ�_i;�n�|�h��̥�g=�W�x�������?�c�z�6a�:�_����ǖZ&��������/'� ]�^�erxN�{��]����T��}��\�(�|���=���7?��O?ΦM;Ȟ\����RC�\IY���Ǘ��J��ne�Q���������W��ei�z��
0�q�o���P��c���|�*������n��[���e��N��i�2����W�uk�8�j�v;�Գ|1�0�pH�R"���p�͋�uHn�{��_zM� ��Xi	q�X7����f�����5(�u�����1߯��S-�\�߲v���������<�����pNJ����MʩSژ�+�.;�����I9�a�6�{�I�>{����w)ɐDټ�U��K/y}=�����Ɗ'�+�6��|���n�Gp�Z��~����I'e3���_,FLeϜ��Wm����M�ի��f���_J���E��v�?s���,^����1hޅdls��9�=퓵��{���Gl�d��J���l��2��l����D��Sy��9`�W������ۼ�^��=1�E�VOU�X�Q���5k��0��;��]w��G�@ H�h�1~�����2�u����kd��x&�M[�0k^e���f���_.Yy��6�[e��[-�*:���s�?r��-D�0\2m�s��	��t6���W��	���h5�8zF���ڹ��m��]ٓƯ��4���>X���Ϗ|�#^�{�f{�ޟ�ԩ6m�[�&��j�O����-yb��Kۺ��N9�l{�%o�l��Ճ[�n��>�4���E��,DԠA��Mo�y�βJy�V>��OD��MV*S�+0qZ���wز�k�З���>��?�~*�+�-�_ř ~������淿e+V�p�W�Iu}�Q$������ZV�B��~�8�$�U�V�+ئ묷��&�3��]��fB�$J?�Pޡ��Z13�fqdh&di���o�����%K<)ʅ_�#@�Q(�(�W�J�ñ?�[��Ź������bG�9m5��F���gj�fգֻs����PiЊ��z��T���A{b�S�}G�]~����G[�����.[t�b����w8���uj��L�,X�B��n,��90�9�ܳ��^�5��|�=����z�2��-���UB�g&�����)���'�EA��?��?{B��_u>N?�tC`Q@��G> I:J�V���D�rm�6>��`��M��@M���ζro��};mݺ5�ӽ���L(�P){�j)�����[��pJ�lαϵ�3�r�fk׬�k���_�[�t���bv�m��b��GV/����|x��.��"O�BK��Q��i��fW\q���u[G�h+�z���1��3��8M^x���6ڑGg��=զr�z������
�Й�f+���)��Ќ�'kNN �-o~��ܼi��rY{쑇��?�gO=�ܵ
�M�2ɘ�SO9�;�X�0�5��~����U�a��kQ��E/z�O>���'�}�l��yZr�&ܳrW�?���bT�=���-��sfϱt��e��n�s��8��R&�v�5ۤ�����̆�;x�t���ٯ}��v����Kg3^<n,���Rv�BV�s�ᇻ�O�{��6n��A������ܕ<W�pL)���~�I��mp�����>۰a��{P�3���Km�aG��I[:�����{��7%� ���?}��?? ��/X�`qw���f௸{�e�v�An��>���b�y�F۸q�k�8c �9�g۔��Z���Jռ�%}�"����,t9�X8,~QM��n�A	 -�����Q���C�G`�G@>	��؇h��K�������i���JRO�`;��7�{�dC� ��syotB��2Q.y,�P^Y �[��f/��#�K}�TЯ�kO��
@�Wƾ�J���[.���'٤�]6��ok֭��[6Y�@�G;utu�o����������sg��46l�d]��R�|���h�\CA&�:�d�⬁�g�,jF�Y���-W�w�������ކ��rI�Z�B�������� �-��1�ݻǘ3~�d�� �>�F8�N�T��x~��E���?OS~� ���b3�\����/��k륤�m��nr�q��#y@�=��I�1��:�����_o(٠�`a�D!,:)�X�0V8f����^!����S�W��6�Z�����Qb�4y�$��N=��<�v&v��8�H�K9�t���v�]��D-R�	��#mGf��'���\n��Vw��!��}����kk����
�=K���c���n��ִ�Ls]V��U-nըf.O�2��}��| ��<��$d�f|o��q�!��)��B�k���.�GA��=��c}c��@_g�	�N������>˻{�96i�D�˱��W�xwa�=��?�w�����������颜�E��¥M����E��rJ=`�Qga@�I'�d�6+D��.e�n�:{rٓ�uTke?��^����|���������Iǜ�$���/}�^�{�g�������Ox�F�9�:�Gh݇it�x6g>��TÊgv�(�\:X��%}�^a�����pކ���z�*�M��aһ���b�Ja�h�T椌QK�ݶ���H��[n���<x(�SԮe��1Ӟw�q�QC���ֺ����I��� ��Z2��g����i��l���-�wh�B�K,��*�)$ӏl���W�&Y�.���+�K�I}�At!�$�aʱxT/����Z�*?�7���l���z��T���(?�o�G���V�F:sU)��M��Ϯ�<�(����@��Thv��tٓ���t���l�T�Mq�q����.��K�ѽ���5�y�G��H>�},���>V�s�\.o�	���A�� 4h3h����i�jq����=P��Z:|ہԮK��z�g6U�V�d�0� h�w�����/�ܣ}p�7 �_i�m��6����ydA�:_�$��03�}g��3�v���iQw��=I�zvvҌCᇲ�d;�c��c͓�"q"���n~������s�]H ����[�s��J�(t����9��\�<��Q�~���Iڵ��8nMg��Ww�ۃ P���H����8�"N<k��W�pfL��������t�v+��N�'�^h�� ��&�|�6�I�Rr����gqxƐ���
�5{�Z� ���\(t_Ҍ�i�hw�4�H�HׂD�F8�QC&#�i�${�(Xh�p��?�� Q�8mt9��=��,�F�R`���H��I{�������ꫪY9�Te3N}%�qR��"����ZXm ��3�;�Y�A�|b*�N4�D(Ś����8b%^+í��÷��0�`�?���`j�T�H��r+�|>�A3ޟ���1���F��q���u�b�|��i�E���@0r�E�m$�4�a]�8Gxb�oT6C�]��� ���[
݅�5�Ȭ�al0����ݵ�P�C��&l܀lB�b��y� H�ูs��_����G� ��|����ځ7k'��c�s4�����"��H���6����|�p�5J���F4��Q	u��Fo��s.s&
A׌��Aɛ	��g���]@0))�b ` 2����
�9K~�z�9=����]�曗@������/З(��I�S�%
�5��`sW���� ܓ�I�fb	Z=�����@���v�q�Ջ�)��y���k��U[�8�!�����hB� ��ڰ�$4^��a��*��:̀?~�x�Ŗ � ����b���;��š�qmX����M.����7��4���f�Цiw��o�}sd��j�Q������
i�~�H#��$:�g?��Gy��G�^"�D�i�wը?잼a;���w���e/�g!_I��Hӗ��"�#����<)%Nt�~��H���zaTJ��y�4�yXL�7n��S)XJ�ЇW�SFN-�^EK�okĺ�?�,�?��<h)��g�����������w A�5�@2v�{�����o���/�0��X��'�ä�$d��7"rX�h�Тb��Do5�rI�m#!�nc����O�n�d~�k��'y�]v��#�S����6��V~g�5�׽��노诊3��)ϭ�h�Q	�=��9</�Bx
��1S?��K.q ��C�(nY<�֦�T�?�C���~�v�d����� �IɆ䨘�ј��\���`l�I�fi��.�b�^`� Ƣpȕ�В5m�����beLc������0eLe0�g��Ɋњt��,��c�. | �u���8�9o�[���mh�с�������<�MT&�DX�p�C�x���x�Bk�)�����8�+�h�l��*i�!��NDD&�z�}����uɌ���{�J���ҾΫ��"(ش*�G�Y1���ַz��O��]�W`�����2�5XK��r������}�c@V)���F��H0��#Ǣ4} ��������=w�W�����Dah/����� �m;��Ԧ������O��ݿ�m�C��<�( ͵�K��i`}�=��z���X��t`�f�i$�W)_	�0t)��`ķ���8��bǵs����G��kk��%��1	!�D��eq�~� �`���h	���e4�M8���&�o|�;��m5L��Ip�o��q��(�y��۳�c�����$+�ͩ�
�CV�Ýު��/j.Q�Ma�d�V8����g+A�O������$�(,Z
�9Gq墴(6ȹ|�(�z�?���τE�j�b��-�,}�CH'�a�/8�����]�v��X�$�R�4��ź��[5�J2�+��#h_+Z,�V1��E�P�%��1pBkС=�C�sW�u'n�^
�<��$�HB���{��>M�R���Q�X�������^�W,�i����6|aW*aMS-����r�4�7���A,�4��c�\s�5u��V-$�<�?��@S���Vϱ��٘�?�,�GqB�G�d��%4��[h�1u�9n��G�ٷ�v�����_����Ų t�	�(�9�:�/�_>Ɓ�~��փ�����pD����빗Ʈ�4���@K��%��"��=�&9!�z�g���0Q���[o[;	����FzW������*9���`Q��^ba*�w�Iiq�I��	��  ��
H�s�o8����U��g��[-�z�q�V^�_�G1!Lrp&��X,{�	���PC��s��`��g��!�h��ڀ7�i;N]����5r˼����'��x�R��OPS����$υ���UO9���M�vϾ���%�{wzI]4���6&sR.���&��8i�Gċ4�Gy�#4H�{����2̳��4ƌ=��C��/}���������;�0w6�p�����w(,E��x��~|��O���1�� bE��p8�'��P@x'~g=b!���3���|���e;�Ph���)�(;�	�q$�F�_L�2�ڇ��~��J��E�J�c�j�;�9�5�����go����6���˓!\�s"Z����!<�����۔t&Ҋ�r�'"FJ�PցZ>C�%Ky"FH� ���&�����L�R�Y4L;͢FHk�f�x�21�)���SO�%�i���������/: �>�E�
`����6I�wؗߏ�1���	E�0?�6m�wN�]xw
�Q�	�j ��Z][��\@IQG
���s����������w��T<�a�5G=V���U�6�d<��z?E��"��(�����d��iR���Md��L�X 9���=���Xʖnų�7�F�  �<Y�R��(Q��bv}�Iu�l�f�:��BL���'����o�g�e�j5/���nj|@��k.�vO��&-.��Ҩj� ɏ�3�K1�9&d�i;�?�6W� k�5��/X
C#BD=V�XQ)--J�G~i.֕�;@qJh���Q@��&����m���x��Jh|d%p<�+�z#��kd�����w�6w��	�JCܟ�'���?��d]�����|�󰁪0K�ħA�1Q��X�_@��KE1�5[�����+SV�q�s�����$�+P��8���z&t�_U69�DU�a�Y��,+1�z6����`A��C(���<�1Yj��O��u��'�d�7���}VhKz����P�֮]��@��t��%���'�����5��o
=�5���i	�_u���PaS)��c�����;;;|a �;�&�@ ��O}�S����|w���b�V%�BT�P�0єp��PBVB+�'II���Ɛ��p*�P���'@�;�/Ĵ�H���Q��9�Je�����@,����yVE^�&y6Y~Ҋc�E`]�I4W��8=UW�x����@�gx뾚�v�'ZNjY�. �!�MTǒ3��;�·R�>����{��)Q]�J�:���	?D{��V,���yq�c˹����c�'�k^=�GN=h�K�^��z>�jmE��AQ!/��$�9�Ƹ؆�@�?p{�.\��B����?]S���>�>t�,��9ȗJ�t*�<hK��o����cB1�f�~�kV,g-�MIF/�a����;�vXDT�r�Lf���|:�쳝n�)�8	�j����P)8Y耇��:�
�m�}�}+���%s�<� R�x%�(>����Gs]=�"������tc���6lp��:{�E+��*���=���q'�^�0)p�gfM���;�Qk�[`C�a�H���`1T��o�����$��������;�$K
��X��O�AEO|K��z�~����y�B�}	ʕ�=���x��9a�u��N���s����~��۶�p��k���7
=�l��Z�ڏ9�h���WY��édS�`۶l�%K���֯[W�+���	�og�=Ϟs�qf�഑FF	g&P ?^��� ��b�U&??L_��|��\�S%P��]W��fϱ*���<�Ѱ1���}wa�h��� پ8���Kt�������AQ�SY2�c-V���~��� �.�v7cރ�NxQ]{��㋢Ě�'A���)�/F��ͧ?��\P��}R�.�)'i;�G�]T�:��3�K�����T�Q�W��(�/�fmA�~������;v�w�̛7�#���k/��^z���O^lV�X&]�'�\b�V���Զwo��`����{��v�igء�fCŲA��w�u���e���.���Pxw3�VC�c�:ʮ|߻�R�l�҂%[�~����{<�'�	�#^,��P���*6�������rV�~�eJ��� Ŏ?�|(�a���.�Q���h�8�����Ƅ;��,�����Ak��׿�NQ�nc��o��h�_c�@��;�ck�x�V�_�-�-V������>h�$�)}op�Ҁ�����:'%p@\8��'�Ē��西�ۿUVk���4x9dꣵ�e��4*ψ����x�b����ݲ�#��+�^�w�(B����A䟀�j��Wi s��W;ː��l������ۭT���N�J�N����vX��������3gz�2�/}�Z�0��8�7�\�](�yS�'ڬ�=�������:�+���G�\�f[6��m۶��Ѐ���&��d�;z�ڂd    IDAT��3`���]����ɇ�����!M�@&��w��Zil���\��_���9�D�Q�5
�=tl� #4�$q���}Ќ�Iʂ�F�_ ���}����[�h7���z?�񖦪��
9m�c�pH8�.ມ}�M�7�_�'
��E�ٗ���z�s;p��g��1s�L����.�3}b_M;k�s��wQ/�۟�2�4j|"������]���wgw�}�7jU*�? �/�B(�.������3U+�6ԷնlXc+V.��[^�D��l6o����y�����\iO��x?�������:���]��bw���f�_K��G�9�>�����@�M����n��.��� ֮Ya۷o�\��:�]�u�[�n�Y���o��N8Ů��
7�]�Z _� my�ƍ��H�yի^� �{*zB��g����*}��z�ȗ�ǚd��T_ ��
�����w6 �Ɔ��;���X�o��}H����w�+�BY�� T�h��rG]+����D�z�Nq��G?�dAU�P�E��u��FT�	�ڇ��Z��������o�AH�r=�&��g��%�g̘�5���|ͺ#T�dAA��X8c)��	��ՙ�O-�AC#�3FPP#3���07�&NX4&�q����d"b"Q.	J�F�^�`��@7�s1�xM��#q�Q�iA��޻����WOq(��k�jY���t�W_���<��>�rP�x�Y��M�Jc�����׭5~�ayy�ik��wW�o�˫͇��7�1�w�W�A���u�Ŏ-M(�i��H���<d��u�d���_�5eʯb��݂?�燆�������M7�p�|���<������Gc�MC�G��9f7L4Ti6|LPg�Ix�f����QGO�- ?�E����8Ё�<�P54 {��G��ի�Xx��J��^fF
�;�?��?}�o���Z~����[���Y�%��:�d�fu䘳>p���� T�8w�~0J.@�9h"�S���"X�6�M�EO�%
ȋ�"@1q���yꩧl �@u��$��3 ��/�Iu<=�("��RC����0�a'ث.��0����7W��>5f}çf�A�������~����ֽo�����bQ[�ߚ:��-��K��<�Lq���/2ш1�]e�������cL<�l>��cӴe�Ow�+LӖ6��ǟ����yo�f3��/��.���0l*�@J����ۇKI:"`y��[-=|�p3c������8���,m�S���R�A�C�台�.����JM7�dG���k]�G����g&���M�TI!�"�'��-�.�5� _un��<
q�|�X�d���Y� �|����_wQ>�f+�y�ր{��,��^ u��M56����9r�5 �V���QG�6���}�|P�.�$a�zM�ii��-M���%n~>w����kk���^�j���g[�IS&��m�$�����u�Af楗������d=�����<�$����47��`h(j�������ΐ���Ō8� ��N��\s�]t4�ܹs-/�;L�>�Eê��&��c�)�:@P����\௳ v�
�l�����MK��ϢH*��1��m%�FA�����V����hH��	2�~�Q�Z]Z��a�����~��t���C�˳᧒8�X��2y�9�G���;{Z�s4�C��|��]��3G�=���>f�wM{'����6�xȼ������N�HF̜��7Ѳ*Ӵ��zZ�Ye�?��UԖ��)S��/��P���G�0�~t�ikm6}*#�ŏ��i���f��LssS�(��ټ��ԯ�Ĵ�yf]}�w�?��*�}p�(��h��1cl��,����F�0dlD5�Rj�
Tz�i�/ �2�0Ȳ
��eec�0d|�,l
�y���}7�ߵ����Oh��;��Ϻ�R1�}�]̅hy�<X�Z��]@6S�Em�C`��N��@_���&�y�1��c�W��۾� ����Ƽ��-�67��_z�x�P3`@�z�*�mNUl�������۫L$��l�3�c�8�_L�>5�ݕ������?>h��/Z�����s�zZΟl�2���!f�W�f�;oϴ����+�j'�j~Sf������6��Έ9���e��T�e~'�kN�'5��xW�/]��*e(��\bU"��r��)p.���
��B�jN=�T�{饗� ����L�w�cU�?�%��^��N�F���_)��.\h���gk���m�R5�Kɳu��s���=7���+��Wz-s��o��k;v��������%ւR�<���iv��u��0��m:y[{��:&u6���'����]mZ[�滧�iFr����k���^��C�t�a�Ǉ|Amm�}E���LY�5����������ϛ��C�d�;[�����7�3ﾻ�������ܞ����io��ƦN3쀃�q�Oܦ/��Y��<��ݨT2rF���*
c��	E--�=��rnfDO�?�������W���(��{l�Z��(�02
�10 #
��5R�]�$'I����V ��G�=���v?`��;Nl���nO�
	��||,g/�g���b��b?ślX��Gٲ�Q�jAk
2���V�����u+͇~`�;�MUE�54�imQ��xɈY���f���jL��l�����y����r����Wjݱ�/Z�h�=���'?�;3�Ӷ��:�/�O7t�����g>��`ֽ�����?���z��N�
E��Qc̸/kF|�M�b��T����c�*Iכ�'k%�e �/!S��Z�͛2�}��kv����g`������m����ݢ�l��a�_Q�����R��B�?�F~?Z.�>���2(���X��(Y�
����qXQo��,�G��œ��>���Q����I��)�FԨj3x�D���7&�n�Z���_�����^5��wXs��:ZU��|��c��8ҔU��:���j���{MWW�Z���2h�E���w#�?�;=��O"x�3<�\p�~��6SQI5/�.v���&[�a��>��4π�M(L�0����8}6���S�G)�Hq#�p�|�@_���������y���!�s��P�}uV��J�T���ϗk����@���J�
HRTUc^�o	��S��8ܞ��M��U6�/�`S�|jW@}��/��v����Z,0�o2�ԟ����~ �?cٝW�-�L�K��U� P*R�M`�ޢ�T$�B55�S���Y�<� ˥I�$ݓ�l�w�3��N22��0~"}er��*󅹄��ء�m�Y�V�N���$9=�Z!�x��}��+�@�t��d��P晲s�ռ��u��4�4���I���|����oжй7�p�Ut�r�<yW�T�Ϝ��Czx�J:��x|���wW���B!�|�!>������U���o[ϊq�zy��4x��ŋ�Ut�����EA�Sy����T��iXm~��L�l(����k�͙��A8�� nZҲxO?���JQlmb��ֳ��ci۾(�d� o] +��o�l�w�y�n82����¸d�Ӧ�	 �߷��4�8Nm>�	��N�� �%����Lj��	��1Gw��{��ލ��� ��\�YʖM+�W��������)���.��gP(l�p�m�ؼiQ��ś3^��s�̖R��e� �|�?���i�(i�.G
�"< [�3�Ea�1�ָ [���@V�1'F�t�_����A��}��-��J�=�5/R��Q�F�8cE��9��T�=k��>�2{Q���x����I��}��r�`/
��!7_2�Z�Ƚ�KH'�I	�=��y�P��u��9)e>�{)л��@3n�eW���d{y^29dА鵵�w�O�2��Xl�iYi���^r�%i�P���2�u��p�b&GY�dA�B#+��E>���m M�g!N���D�p_���{�9��]ֆ�g����V��:�'VY���o��;����,O&���%o�k��l[��WXA����[o5����=�@�a	o��
�@���)�٤,X'Z:c�1mf��OA-Oϥ6���U�/`�����R����n�=2!0���f������<�J����?� �?�ܒ��u?���+��s<2���;��sm!# i��3�5���� BN~5�����IgO������H����)����d�k�0�k���y�f���4L�N�b-�Ħlz~�Y޶�8�:s�J�3g���@>���yF}�����K?��/�j`
Ɣ��xd���<�U��~;>�	�i��HnZ�<d����u�.>�8��b����2�m(ֵ�N�,~iu*��,"`ON?�}�m,hr�9T�ŕe�=%�,�[\"�c��h6n1�Bl*�q��������m2��ҳO�4�o斲�mO��
�;u
����S�>m��WUT����y��l&)-�k���x��h���r�=�	�]*�g����q����7�^��\��Qq��ѥ�v�`�x��z�H�\����SbN @��w_R�Re�} 2d�,�=�.�(�~���chqrޙg��>7Z�>K\�b�-�1�Ϥ�d���[6����c2��s�O��g��{}{�F)ɪ�QCCq*#@ԩ�J~b����w�� pƃGKJ7��Fź�]�}������C�e
Ƙ3)>�xP d��ٯ(�[/Y���d�Ew�O��(��N6�P��&�_ZWՋ�����4��>�$��92a ���
S�xJ���j�An�� (
E�k�IG�*j�T	cM ���u���J�rS0ڂN"nA�GQ����d|x"<'9�|�R۸�@UHV��R�6������*�Y��&��
�G�bL��8����]�Ck!��뤸v%��'�LjL�����di�&s�����҆��|����7�W<+� ���E7OR}�1�wJpd� �6m���3-��d	���'�p���/Y�ʣWF�֒�g�jf(�M��?8��,���3�z�V�T�2�}O��`��KT{�q�x�������^a_��`�^c�6U��Ŀ�E�fƈh_�oK��simm����)S�b��og�d�Xx-� �u�]Nյ�e�sf�YH�G��ʱT����D\�xg�ϱ�\���?��u��a{k��`|?���|��M���?�����pc��bG/rL���	@]�������������B���y�~ �>�:[�L���}{��~}}�H
R���񂠜Di���������"�2t�;�ȋ���Yw����nv����3�N��q���F@F�*��z(}_YW�||�Z��|?^�&t�,X))�����:�w��7X�^s�g��W�j�	䛗xz�${�1��Dɸq %> ��)) "�^Jo������/E��3�%Ydb�0�k֬�^s X�c.�,���7M5)�[ލp@^�"�H{^�\�EJ�>��-�������ű��)��_���@�)��N.g,�ׂi)3A��I�
�[�wJ�k�
tt��o}%ҁ%��r�c9� �Ud,���J�g��R XԎ��x|��tM�����/ZŢ͐���O���>���
��e�5�@���f���l�o���<3|�a�2���gPX��Z�?�Q��8k���ڂ�9����z�QGٸ��5�*��}tϋ҆:ԚBy�(AY��R�2p�K � |�M��K<��ISK����r�
�?�D�7�H�~�<���=��+�����9k��e}\�'��ε��KE�6��c��갺y�|])��xc�l<�ﴷ��(�[�F:��N����b���g~?����Am?s���a�R4�.nHaK!
oDm2���d e�=�Sy�:s�E�*>�2��X�qj6�( ��L����ܝ8�dIZ,�A��U�h)��7�{��J��od�5�CX ���{ �@��թB.m�*�Y?�ļ���nu8d�w6��!!�6c�!��象� �x"����������,}ι��=����$_���e+�U��`3纲A�lN?�ck�[��c���UJ������������V��D� J�C �~D��PV�A�+D`��3Go�����!N|S�f��D��p�}Cn>�$0��(*�/Y�X��/Xʌ᪟α�*'����d��k��"� ���������s.M+c�k�RgϞ�ND`O�	�-ݚ��d^dy���Y9��h<cP���衇ڸ�G���R%�̢.?�Y���\cEϡl#)���Z���amm�m%�O�����d�?�kd �X��d[ @���� ��ȹ��z:��H�:�`�m(��Q�6֩
L ��+Ț�Z6�F��~b���2b�� d_�m�@�����o�_)����Y	xc��I ������Y�� .:��� i��Rb�����X۠5b�?�я�gB�(
O)�xU�.2$\�����s�A@A2_o��Ft\����͂s<����{sv4��1��O ���� ��/À7��IW՜s��f���|�i^ޡ�͟k�H�C�"�,zf�����]��+Gm�0�JBI
�ˀ�U2��}��naݭ%����_�?V,��SD����
�m�`
�@�2��7����s�)w�7%%e��r�-�2"�!P�����L�����Oa�����?c����k���8�kg���O�1,�Q�F���41"����ǈ@�g��W2�I���\?�D�Ld��Vy�J]���|3>y��_��k�I]�O�N�VLbW���<��kkko):�<e�c�����h�]�0;���Y�JU�u8F\m7G�;�*�{e)�9e��9l�N2��;�;,�s@�Ԁ:Ԅ�����[+?�����9Wm���l��--�������Y��?��mV�G����W�})�".!�������H$}�D�'N�'�W���qO�X�7_�����}�`�h���В{����ߕG)�P�W4����7{��1�}�����̪[�h^с����o�&���O6�w�'PKJ��q�A����L�/ik��A�?�?����4���	 �^�������F��ˣ�>�\q���anPrk 7���	����s 	����K\5��B�?�r.�$�W@� .� �,(�ݦ8�b>�d�'{�TfёPrx-J��	�fƸ�3;�������\�����(�Cr,��Y`C�� ��|Emm��%���h,#,������
*+�$|�ff�*���m"~�}6ΟTO����(`� �7�'=��C���( ���PN��p}��e��{���x��,��Iٜ�����?�NcA2�|i��Q`�!��CB�3$艵��@�9c ނ|)��A�}��'�M�m(EdIVv�\��v�.���)��w.�_��x�����(h+�'S��d���Ʒ�ͮ[TwS�P��g��ם���5bQ��[���& ˆ<���m��
oد���dc 초����-��!(�!Ç��j��T;2������g�W|�8X�>A�6�_�	�����	Z�fX��z
w&�KcA�'���R�$�
���^
��"�f��W�&�C��^�_5��,�w7#&׶앩���Q�x��񳁿��w����*~W��(�ނ����S&�6�b�?�>�( ��<k,,�P�Kr	�6�r�*/I%�|h@��*<�N�Y4�8)u�M��1��M)\+�%��_�J������@�o	�}P͕��Z��1!�MX���?��r}֚���Ɂ�'�/y�Q�ɋ葇ӅK�c�C�4oi��#d�'�T�jŐK��ݲ�1n�I�t-�\��˂��*�E��mo�zO�[��?)��CO'qw��;�_�� �y��6���m�6�v���KdEʢ=��al����w��%ݓ� R���,.�
K���'e����w�%�{˟N<�B�?�?���rD$�Z6`���`i�    IDAT\j�'���@J������@ܢC��1��P.j{�ߩ ���s�1��d\1 ��y�.��<���������ɤx��D9�j�He��.R�ʣ���Ӥ��Naw��z"�-j���w�9��������:X�8�^X�p��9V/	�@��ķ�M��|�K/1���;����{��M/��\�2>�_U��L����](	��9�\h���� ���-rÒ�(K=d ���v��W^wwy�=ɔ���{s����3�.�e���R��t% ����yE:F$��y���/���x��������Yg���/�˳�7z�@^:�2���q�SEn�<�WM�,�'�|�ƕtɹ
����E�6��M�8hGɂ����ރ�Ҹ�]�]�y:�2��E�a���)Si�5��
�_@Z՗�'mjDux�(�Bȱ�iŠ�Mq��բ@-�y^ �9�?�n @W]lF5�S/��x�0��òǺc,�r+���/@�kh� �����k��w�A�(z������]EQ��/pI�d�駯yU]�LGb.s�*	? �,B㩫+S��52R
�x�z�W��ǖ&t[0p=�} i��B�P(�G� �T�r����}������9�w�F��Y�ъ�zRT�5j�o�(V�+<���0��������ŗ�?iꔇb����S�?̓��`�=A���b8u�+��T� -B(���-��O��=��-<?����<��s����K��d�;�?@��/}Ɏ�!��q�3�=\P��ML�7���;�$�K��d{�m�l3CRV?���~�^
@�� ��?�{���ώ�K�S�bs.P�okB�/T~r�F��5u���]d/�~��;�3�?��24ħ�� �mj��R.R&:�:�X{C�=�<��C:]L��n :��>�߿�GO=�D�w�<e��i�5�!��)��V:�
P#����\RH���XHV���Xx+V�H��U.����	����`s2ר���sp�ƹV�I�5���a�A?���h�"[�K��P��#&o;�KV��)���y��S#�<��؊����c�  (�����l�[)��v�gw����u+b}�I����#�ܐMƩy��� pU��|'ʜ@$4�:X� ��c� �(2��3BYI�!P=('��w����'�H�v,͚�{f���O8�������ŏ_?��S���5�Â��v-��@3�� K)�XH_��K��B��*vt�M��f`#�7���j�q�]�p �i)�����e~^�� Y]�8��a�Gi�P3:>�s��w[AwG��T�BQ���Z���P�� �m%�_�M���m1^x�U��T��ۄK�/V�w���a�J�����j�u��\�C����:~�Oz����O�|�^ �뮻μ����j��?��F���;ڲ��i�9�5�a�o�
���{�N�U����S���"�V9D�v���1"`|]��;����g^�0����|�]����O�')�vO��Y���*�d#�	A�{6  Ϧ@�-�ʝW{�̞��VIc.h"��s�Il:�uF0o���ҍ�Ld|6^p�9���`vu���#��5bx'��k�eA��I!�݄�/��T��\p�����r� P���S
�>�\|�V�*O9h� ����i���h g.�I�k�	�gm����?�Mx�4�|��Nu�d�-|��U�(/Q�Ɍb���.����j�����l=����x�s��a>�У�)B�r[cc�=�~XX�x(����mm����aWf�,���7��T<�VV�{������8�b���ӛU�� ���X��lB62uӗꇱ1F�1��6�!���(*p��#�1�?���R��ݼ��<��)N�˟��g�.���,D�e<sQ�r��$)�C�s���{�N�H .OS�G� �oϝG�U���2��N[)-Q4���߅|�{d\j�#ߜ ����I���]9�U.�x�u���u���o\��-���L�n��ƫ�T�OgJD�v#!�X�X�:��M�S>����tK7��0!��'���@�?�B}�y��C۸��5�Rg�jL��;����+} �j����Ac�Z�j�Z�|k8���-�K��6P1�?����0?�?��%�-M����8�Y2&o��e��d��1l|��	��t�WkKO(*�m�>�g�)��ؖ�Ke~rO�_^��+Y��TRyԒa�0�H���>���[����4�/N�k��������oO���'�3m~��!�m����K��4�":(�'V��$]�]s�VѲ�]�K�#��Apw�M��`���i� ��z��d��]#���Wq�֦n��.�W'11�dz�y��f,�yF2MHC$3��J|�Q�TO8��LJ�J�eZ�C�馛�x�����9Y��b1�7�с�2����x~h}WZv�er�g�X�(`e6�5�<gbܬ��;���^����w���a��3>,h�V�#{���O�~���z477x�7�y�O��7��Ͽ���^_������W���Now�Vs���Pv9V�<��5�  ��'A`0��O�P��݁��YY��=�!��( �� :�Qx(�8������K'�i��o(�e��pjn~
��W�=�%����g��y���`���yꮲ�>��������ᕒ�C\�s�Y���1�8Lf�ܹ�������J����&g��w�1�ͳ�<�[�w�ڢ��|�G|������l����=��]s�����ٰ�e���8d�����)k$},A>� �H��f\46Sa�t��`�ɂE�͘1���~hSr�� ]�E�qh�[Z2�0�^,h�rt=�B �����O�Q����k��?���y�I�ĲG��ƿ�� �W���Jnh��}d��k�i�X�6��mW�|D%�g�d˟uW�+��θ
����e7Ͻi�	�����9��˗G������۾� ��"���D覻;�+�(>�wQ�*+Y@'�7����lyv���H�� �A"*�`����)� ���;��������aEqo
��P��>H�$�"CF']1&�
�����߰�I���u�.�ÒgO�g.)�c�PH�A� J���w������$���o[o�އ�=�3c`Ȏ��x����.Yzaw���3��(��O�x����Y��P�]*�W��-vw�����С�d`(8���Im(�_�)$��͟6	��un��RN����c����= +�-���q= �L��Y�����KA�����Һ@ֿ{���f���8ԅ�o>�Y�FoZy�V�?��5'�S�H����'D�
�WZ�^$��?xg0g�l��T�2��ֶ�	��y��=[���5׌[��s�Ps�ҽ2b�Ӽk����_i�n_ײW���b�\|�S�gf]�gm<�,�Ϳ��J������a�Pm�p�B[��D�?ܿ2F\�E�|ƯϺq(� �5k�=xE�\�	TP,��]/��C� ߮'�{*� F��d�`TA��8���6̤%sp
��<M� 
��ۓ�}���7��Omʭd��.���rS�Y����7/�q�)�?㌕E�<��c�}��~S�J@���}������XG��4Qt�jS��|�3��<7cb������%�����8M�Hl,��*�����Z��w?�Z�����d4�����¤/�I��yEQ��"Њ�̳g�>n�:�Qv��?�?@��!������Vz+nB�k����ϧ� 뎼�P9���s�I���7��������@��ͦ�~e2�s��o�{�-�A�����ڴ����sX��R?p�z0ϻ����`��"q`!���Q
�R�5�LlO���SdD�/Y�
�a	`j��P�?�x�Ny������#e��w�ːB�'=� N]�tU~RYK���eZ�x����?�wPH�h���T�>�ޟ������/c�R�������<��axfd<�_�}��˵����q��յ�k��o�qyу]]ݨy��-����6 �pQa��%`^�޽�孱���&��f���t?F!�k�Me͕5!J�9���LOr������ٹs*��wS%L(�2Zb�����9p�pǀ����Q$V>Y.��
��J �'#��cUc�B��=�>3�a�ųJy���ݺ㡭6�N��3�����g�bW�G0n(�y�7Y���(�"�L�//]�9�O������~H��+
�2x�Iz~�p(l�xZV����]�.�P�����z����s���:l��t��m�1�c}Y+�*�tXŠhT�{dUQ�-���lsR����~�UH�b�T�j�\�ϧ�rʧE�L��i��[�z���x|�N��F�
���%m.ޚ�G>7�c[��[����'�! �r����>N�K�\��75nN��"�)�&�w7�����E_��<U�r����`�*A�� ����'U�X�|�@������J�T1���Bʏ;ܟ�S��HhO���<�h�J_Ei��g�� �')�/���y�駶i얹�p�s�J����!�#wj�)t7��w����m�������-P�ޙ����
��a_�l��+��<3
�y�M���O���ȅ��HH(�\tw/��XEvvvn3f��{��/Z��*ڇ�_�`�~,�;O?Myy�; ��E�v �F�:�r�7�Y��>xܸq铓�LP�tEU��˃E(�Q��m�UQ����L�|��L�cu,_�Zuڤrְq�f���yq���.��Kyq/�	J�MN����g�B�j�\/���t��m�V�*\h�p-v<z�C��l�%p銟0^�}��Ȋ<��s��3�ِE��SOn���sJ�?��/�0�̧*�W�[�gf�Y�&��-CF5̽���ho�b�ʬ� ����q �]�_�N�S+y��DQzmy?��dXN���k�O���O<����\~��ǿ��˿�ӧ�H{�meEZ�܉��s7C!�����r]^�,0�!��e�a�;6����Ea��Wm~��_Z^V�"�Ue~[]������TAO�M�>��yYm���㓲�d]���D҂?�̼(��!&`ѽ�,�^�	�wQI���O��z�(p͸�QQ�'��L)@�O�QAA�>���m�E�06�g���4ߋB�Y�lN�G�b�#c(��z����`�R�G"w�� \zO�\4�s_��%���}�q M���p����_��| �����U�<���^ߵG��Rm���rV�?��y���)h�����'�|mCC�%����9�J�]��K�4��D�ȍg��:�hk7��~�3fL�e�F�eVL������}��g-��� ��<w�)�9(gS��~7��sdZ��m9� ~�6(�Ϻs$��C�v@�����/����(%'�r�H
Yi�Fۙ�5'|ʊ�'2�zi���~P|tO�z�q+;H�,E!X�����/�} 8r�a3�%�Sͭ�S���_~W�T��p�G4��h+���kC���[�-m��ȋ�^d8�.�K+|ݏ�j��.�3k�Y}�n�<�ӯ_����_��#��ܓ�/:�gRx��!,��L&OE�宥�����=Y�\׈��e��a�6iA;��@����<����"j�,�_֢��I�ϊ?tw��y^�Τ�D{$y��M��pĔWT��]��d�+����w�G���a�1?�ݑ�v�$4�X�:V��x�_P�T�P��QO(��K�R>��9�oX�dĐ+O!�㓬��c�+ݏϋ�p��֓�c�/Y�����z��B!�G&�%=�C�א	��UUU՞�<���:
U$*�=�]�s!kY�e\娹Ҙdd�������s�(�C{j,'�A���sT4/��Mw�W �L�%��m�ng�J�gȶB����%���W]u�'N���^E	�����_?lٲe�&���P(�E�Z(�mƠ	-��|�����
�d��
���cҜp�rQv|7����wb���-mQ%����/@K��*+��s�Y�9bd,�G:;;�^�y�U�!Qc�6lذ���/ZB����,:ml�'�S�G@�^�������ŊP��6Q^����B���M�Pn4�#�5BqṸ���nZ�ƪ{�l+V�X���}�z��6TVVvvvv&����x�kkk�.qsss��7�<�����D"1�ϩ�R%N6�;ǢQXGY����E\/%�idz�?��}�dp���ʢ��mŕ	'�Tb���;]z����P�+���TC�ВiӦM?������E�L��W_}����vk8��#�b�Kg�t�����u��7+@R���h�vԑ㶩���=l e�P����Ӡi���.g�qh=C�����)P�(-��O���֯|�+����y���jmm}���	�*|r=9�f\�R:.5���)��,���<{�g]�s)և�9����Ҧ1�J�m��u��ׯ���c��3��,Y����n�<�L^TQQ1P��F@�m�P�R)))�LP����nR>�����^����I��C�6�#�S��{K���!X��V����>�Ogg��&M�����/;r��&j�̙_x��7~���|Ruuu9�� �+���L�uG&�7�u9J崓�uhS#c�y�\�6 ƺéM���V�����ZX�x�O��o��/�~�ĉ�͛�yPvwwvv� q�xpV�y�mv�����92
`� `}}��	&��\���5���/f���\�D�)���K�i��5k����WJ�QG�{b�����I�V�y���	<>eE�{��vw�()Ŷx^e7��ʮ�3%N#E�꥕����&L��ùs�Ο��H����Y�f�O�YUU%��!(�rPQ��Ke��=hs�|)v�J��pD'%���~6S���
���s�euf~�P��VvGJ�mPS�ȕ����1��a��{�wP"�x���k��/�uQ@o�fv����R�t�u�]���N8aNO���g���[n���h����d�E��Efܽ o*����\��mI5ֳ�AEe��� �:�*���������'��(9A�O*J՛H$:��˞�������:�����&��;o��§gE�E�0�:g��M 4�S���{�.gs(Sg�j�i�e���E�p�����M����8_�?���W�"�HcMM��ٳg_s��Gg��S���1���NS%(��L��<=N8�閿K��A�,׭[��c�=����|�w�q��yvuuUD��#cU��������i�lRY�/���˭�p���|�S�Ac���x�{|�ғrPFolll8p�G'k�܋/�8�>�5��;����O��������G�WS3`BWWW�F\�@�|a�I�m�P�����o.�W.�v  �O�}D�d)��H��~��UJ��Xuu����}͸q��s	��yh�%�+�1�(h+�_ ��"sn ���[���	A�$_��*풿�8��L�0�P(�p�'|����Λ7�Ɩ���*��?Q�W+N�o\HAle�Q���ԙk �2ʌ�� �έ�����O���gd�RJ!������C�wڕ�>sҨ�:�z	����n��sK�~�g�S*+*noo��!J$H��6o>��g�N����~�K�2H[�X��&+����t_��� p"[���i�a��[��kN:餜TOj\�c�<�+̯,~Q?���xBA��~o�_���;>7�@����q��{�8��C�P���:��˗W�r�-��dӧ�VTT�+�\oS
 �s��Bge	+�!��������A�G�ic�{����lR�*ڔկ،�&����k��j���5gΜ���^k�&{�=.���#V�Z������-+UQQQ#�I�-�Lv���l�&�|7�M�e�g8Qy6B��>�΂�$�������o��7��>�z���d2�`8>��� �G֒� ˾'߷'_�&��A/)�mݸq��cǎ�rG-�ǲe����_ߵ���*p��.�+��̜�H  �IDATy�C�T���>��/�V�	$v��Lr��^A�A�	��h9� ��ۦ��������:�����g!���=�͟��g���u���S�x_����D�	�BeA�Y��=����$�t56�/碌��L�l�dM�B����S>�+�r
��M&�=u�W���O��ӹظq�QMMM����k����,)
�h��+(�#�z{���9��3f�V9�1�S�zÆ�ǎ{��X�����ȧ�x<>����wSi��1�}�qf� �A�c.�WO&{-�4�S�D�o���}_�-?m�p�)2%����Æ/=dԨe�_}������%�߁�������y�o�f�ڣ=/1���r0��1������G[_���m�c������X��l-�d�+�F)���(�!zuvt�C�Y��b�!���dk�,GnL(�[�!i4e���I�?o���ow��ߞ����[��0&��x޿W��{�ҥKw(?��������YC��h�H��СC����&�Tjoo�ڰaC���2���E��]�,K�·��gw�}���9C�2g��i�������p+	�{�����[B��F��^nhhxvܸq�������˗W�����4}��}C�P�"��}�z���^YY�d!C���}��uo���߳�dS"��������(e���3{^��8����Ic�e��m7���D"������5;�Õ�}]���m��n���Vw�X���i�<�-�յ%�%�G��F�<��G���СC?�6mZS>k���R��Ʋǽ�dɒ����������6m����N$�
��D8��ɤ�,�3&	A�d�/[�掻�q�{���F��x���a��q@�1i<�Θ4.~2N���O~�߾��"a�ya/�¡d(i��ԘӲ��1&�������pg(jO$M�H���΍w�}�_�������w�jjjD�����Ӳ��pWWW����-�d�-5���ye�%�ɴ��L/0�LF��p��<����T�B!�3�L�<��o��S���z�k����9��K`�����RH3�]��u���d2�Qc�t��y�
��P�q'��L&�{�GH�1���J$�Ϝ�e4jMd��:��h[(�t����9s����px�>}jR�r�|��i��~�`���/o�{����>ӽ_����R�;]�lV�<�8�dKE}��P�}:��%�:]��ʪ_���TD������ͻ��]�0s�ѿ'.�{��k����m�lI�w��Qm���*/-��'X<��j��/�Lߗ�~N�Iw��~u����Q�G֩.�~NU�6t��Fc����q���K<"y���!��ˉ��g2ټ�OJLI[`��j���A����mP�C����X��9�?���cfAt��S�b�b��_)��%��i@k���1O=$���&,� ��~.�� PK   ���X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   6}�X~��k�6 4 /   images/663b53f5-e86a-4272-a51e-f5b809259b46.png�yTS��6D��U0�*�n�4JTP��� ݠТ�
A	CP�y��j��mQ�L�4�@ ����@E� 4$"B� ���пw}�ߟ�ֻ����^<U�k�g?��u��/������[��O$'nE%���W��o��� ~,=󟟏|F�W>𿿦�t����G�ɩ#��/ׇڸ����;�7:D;s���(��_��b�	�3��G"2G))�)	�-�H��[_Ɨ�e|_Ɨ�e|_Ɨ�e|_Ɨ��H�<�/p�������/���2��/���2��/���2��/����bl�9�Ϸ �?��7��S�9gζ���Mт��řv�����'�6~�t�y뽇N�ugKZ����������E?�G�'���O�0^}b�r/��̪�=9�����g4K�?E�d06:�b՚*������2��/���2��/����6�!7������CSoo�Q�ا>�:��3�"�ܾ�yT�_Ƴ��1\�yk8�v~�V�����g���d)N�.�х�I�3L&�}z��U�B����I����Os���:�O�@�bt����j�A��,��YZ�Qr�p��`���5��^Jt�l��3g��g0�������ҀŌ��~~�hcG����a{	|�K� ZZ��,��%�o17�����2`�`�~r�p�*3�������(�w�2"Ɂ���@�hy��ON�����x�*���/lU��b���].�?W�-�H$+
?����%{�1��x�EF��*�2��K����AZ�� ߸�����4@��_0+��r�� ���g��O���D����N�ʲ��\�C����6t2*�vnȺ_`�",������Y�;����Ui-j����L72{=��H�5����CB�:�F;���k*�3{vaa�q5���[X@���n�2T7Nah���-$NTײ�ڐ�����	]�8�scO�*�XwF��)(7�x��xλ��r�	�F��(��s�����1�QP�Ƞ~���4*��M<7p�'��Q�A�����"�t�A���t���#ڇ����l4}����c�v����b�|bTx��DǑ=���M&BI�$������.�k��>Ը|�B���C��VQ	Z���L:gO�]9����C'�K�Q�x��ߵ?^˫�S��ai6Ǘj��:ٗ�`4|x��Ǐ�_�~��*Z�&c'ո����L.����\쓷RE���a���<�g�$ݽ��̈�r�3'�0J�����:=�3#��a+�^�V��65�Lm4�����Ne��w�7S3�9�70^0�͈����Y��K(��34=A�)WB�ێ����%`	c�y��j^�1��!���Rc�	1�'��p�<�M[`L ~��*3���gϞ�~zi�����'��&�\f�1#��4�j����]IG���C�������<^ֹn̎�1;�CvOm4��bD������:����xY9_"�ğ{t{[!��9�	�9�^��I�s7��'�b<IT��V��1 �y��lb�H
�O��ƞٍ�݄(�S@���<H����$��Q���������*�� jA2�Zf9X_c��i/Gӵ�����={6(���������	�#���Tr{��@y�?~�O>����~c/o����J\��ê�Ȼ��sQ�T�&��`j�11�<�C��,��
NW�M��}�*��<�~UhNHLө�����N/M|z�u�~zԳ@��}�<9����>b�F4����eЈ��Ӎ��֧6��0��D�z���j�4 'O��
TL&^rd��z�s��?�iV�c���4˼��i�����^�� w,>�qt=��c�H�����¦�F�������To�z�b�!~ԅN�m��m���NAn�>13��wSEB���H�zE�^`M��F����W +6fo��I(ƽñ�5�!L�~q�"�qP�ܞ̜��g�A��m��+*��-��f����-t�3�B�u�9��`����5����h������;�s�F�,���Ը���3��G_LY�f6 |G�����#��n#�[K�Dp6�x��}�o�=�{��x=��b��r8�r'6�̉������.�\��]��wz�;Ñ��fG��l������mG��C6�$�'��]���drd��ߘ�F�/�M&&�3�/|N�^���7xօP=\�ۭ�
2�hƩ�VS%�w��>t7�ޓ�lu�;���+Qm�YP�����D7y�s^N+/����{G_�\��F����x�|vv6���	e������?lf�J�����ߧ3���_��- �:�~>�fE�Bp�:�|G7ӬEIĕ�@s�&9��ͼ
Q33҃t�b�\v��=��7f��Q�n�C~��^��ӯ`K����4d|c�3�p���2�����|+3���MhN�+v�՝==D恾_��.6��3p	��w�t��(�EE �B V`��Z������-_8��w4ՓL�VJ��gLSɱ�eq�.E/�v.Ϊӛ`j��������]���	A�u�ݾW�jS}RwCu]7/���E##v##��-���x�'w��}M�������r�E|+��Ң�����A�@Ɋ\�Ew�{��]G�p���̙d�a�t��,m�_Ѵ�����������_w�F/�PW0���Idjw/�/��0_:���}��9)�s�
?t���qt:�SS`U�jh�����]��?�ÀBj:�'��/0�����q�<쌮7'Zs��u/�jF�>�U�,�T�;�O��E�t"�qF���o0s(G�FzQ���jpئ�sY�c��'�A��)fNkK*�}���ݶ���ej�W���p:0�
n�I��,��،`T�QR��W^^�>5�9���=��*��U�쩔��mD� �y��z�E)�lA��i��v07��r�m+������X4�;� ��?�ɖZ��הhiSS��%�%X�C,���:\QΏ�$,���.������?�.*�*~XW'�KVw�1���s��C�J���|ud3���F9��{��̈�EZ��B9�If����O���0�O��K�B�W��6Y/�>��X�[���]X�|a�{����x{ژ��~-��b����@W-��z6��
a׾b7A��=m ��g�26����6�K	�bq�H�	D�	��6�dE��=���f��0��܍�!뺺�ɽ�F�������_��Ved�%��<��陙>��"
0v�:b�(Z� �F�����cG 2T�ysA��0-�Z֙�O�U�Db��L]��,�Ί�֫�����J���+B��&��>�e�Y�X����<��s��y�,����r3T����H��ŵ-�ڋ����y���ڨ�eO�Cql��G�a�/cz�f�l������~�����ݻwS�b��,d��n���0Am�:�R 1���L�".?Ƣ����w�j��橐�]������+d��b/�S��E�JlA&R=F]8M*�.�Y?=�}~W��ѣ3��l�t��[ I:_��,���S�NBG��S���Y���"��o�E/ߙ�eJ&��#�1�% �0�t%C��y�n� �G�Z�="��K���LФ����?���;�`:H���pc(J��)�`��bL��ئ�ZW�c(G��`%驲v��j.ڵ��������B��@>���k���\�7�,�h��յA��{\56P�O@Z�'��!�Ȭ�@r{��H
ڷ�K)�!�L�� �;d�f�i#u�M��y?���A-���,���W!��x ��Y��ߤ"Ux[�'(̌�y��Wi�L�DD�u"##�o�R����N���"��&�����?�ݎF�"��p�U�6�E���"%���u�s{}�C��oѳ�A�����踙�7�C8�VO&B=Ȗk�Ҭ��o2�3Jk)�m�k!(�̒Tn��h=K��L�6a�X��Dn��)参��9}���Hr�2�b#"h#���
���Y�bՁ�G�g�uT"���+��Z��U� ?7rX4y������<�vP����u��$�F�ҙ�.�71��
JH����}9 #6�'�@'�tHc�B��Ħ�>:@��xB@��fjY�?A؁��M�ΉN�aY"6W����1N�����=t�����{�Cn4d'Q^���Rۋ�b����Ug�ꔵ����������[�V~���s�1���Z���⩑�S~���'ZZ��+�TFo��O;�pZK�J�$q��Q����U�j�0Ys�I���D�\*sfpp|Z�p�Q��%5Һ�3n���?�Ŝ��{�����n�1;�T���0,Tl�Į���.��oMd��%Q`���ۉ
��빯Gd�FL���=�O��+D������C�y�`��>���D���M65�&ƠV�3��_&g�2����E����A~q�_��j}ʹ�vR(�ܿFP~f�U7w��G��%ݩ�w���J�2]�z��`���-TN�-^=�葆�R��Ϯ�K�7:5Ǧ�58v2/f������\w[f���vl ժ�?+ ��M��U_a��@�y��TF]P�J}��</�o�d�(b�'��Ю�yi��k����t�RI���<x@�bo�w4R�i�z@���t/L,�l��Ż�E��9��#�P$̔�r�����n��D;}6z�:�aC]��r����^�� �ÿ3��:GA���������0p4�A����/>�=OKcv��'Y��>=G��:'XO�}܅y���k02^�-�>�T:�z����~4RN��蚾=�=�x���\��s�����4����ⲟ�u�\kc��e�X��&L�a�_ �[�sl<M�u�yٓ�,�S\��Y�41ܪpk�	ޖ(j�������"ń��>��xG(S<��]$��s���T�؄���o��?���~sÃ�#��= ��E�@�����Қ��b��Ӝtz!b����t!�N����ǟE�ȟNv��������� ��.���ZW]z" 5Z�~i��co��5�b���ͫ�q�y�[	����R���%F�b.�|	9��k/�&.����������Q
�ѧ?1��g}䝍�&̘(R�-i�s����5��W���'���X<��1x��_��'DNM@��tu�u��#�W��a	��������P�34އ�`�'��R��I��!�ꆔ��쓁��t�jl$���"6_k��xqRV`6���l�p��Ю+ Qe� tW˿yr���!�/���'5��c�ׂ�4J� �S��G��#��7�D͑�>���`]o=�,�t�9��=R&�MC/ӭ÷k�rѓglb�jV�Ps7��t��1��rF����A�%\��9:�}����g.>ygo��E���|����n��ٟ�~�QP�4,`	y��7)b�[Jpq���1>��V��,+��w�^�l[�e��,�U!�4�p��l�쪍y�-^y{�9oP�E�f�o���*����͆���|���^���X$�^�e������`M�K�x|,���s�}�Y�T�Z|�~��_.�)�j�̴bī1�E�
zvG������`�\�t���Fz��s6��0b��5��9���~�_o���	���?�h�K��T���k����կ��śĀ`BZ���Ț"��wQl[x���	gM~�T��&�͗�6��[+�	}��&�Հa����0�K��=PP*��0^z�n?����S(���1So5S�Y��E���˜I	��avS蒶��ܓ�/<D�����#�eޙ��
M6$�m'�c��݋9�gw�e^ڧ�:5ma��o������b~v�C�{�W}}����JK�UY�
�Jc�yccc����<U���E���9YL��Ւ���wA�e����Ë=�E�����*	��XY2P) ��-��t)8aKj����ж�*�vk�dS��XZ�@�x�SSr����D��Z���,�x�M�}*;�0p��iqjʥ��o�y1� ��G$#��N�d�zK�2�}(��?�|�u�V9�'A��1B�nG6���kD��c[ݎ��Ps#i�b� W ��->M�,?�'�!�� j�a�[�`�8� B�8��W�/j6��%�C���b���mܟ�:�B{�����������MaA��Cq	�k�
���&h(%p��a��AXR��~dM&�h��uR�������,sٻE�H:
��GDߛ*g:�	�_��[7�&1l��u]�W�2&�MXo�u [ �p����d�Y�C�d>��w2����@+(��T�2�#�@ �)cF�#,0 �^�K���5�j�D"����;U��� Egȏh��}��B�t%}����G��27"�0�(���I%�:�8wGd�fUUպ?���6�8�Js�
��)���-�@�ʟ�G�ز&�~T�C3��^��suc�4�]�ɖ�Ѥ{�"@|3��Q�&�~^o�l����x��%D#Gag��n'�@P
#���u
����b� ?���(���13�~K������6LH^�o���"�Vh��c��?����#5�QNiڧ�NM��JwJ��Z�#�񿃏�7��𨋙����.� �l�=�")ox­�$s�����4�Q�t�0����c(��dJuT/�tCI�Z�kP����my���E7����zz�kC��߀~3��>t�ҩI�� ĸ����T{�z$~�*�z���4ˡ��?�٩�,�w���h�m��B
�����g��]Cc�YT#,�f�L����"�<\b�h�͟�+�5MihWTG�am���E�i���a�B�O:	�˹��y?�dc�a�"�Ƙ�,�����&���d
�Ks�i�@��v!��6�Pq!9T��3�U�U�Y��j���L��2�o�1�ڊ�[z@��������S������lz怒���y�!����������#�v��)�A7��ߓl��[�;=��Dy�d�`����@�W�|�!��a%�H��+ȉ�m�'t��1��0�	4��E�^���l���#̾�ݖ#���yaA+]�ۿ���O����a˶�㫀�ܹ�Ҕ�P���7�U��U�����P6�#w��'J�kC7�a|�Z��XS��A�	:�'�9�*'^<31,��;�NV��2#� t��;O���QpA��%q�'2��<g@�b��G/˴uu�� �]Z<�������
�=|��`]W���l]|{�E�	�V�d+��Uw�r��x6�-��h�����*uтj�j\O4�ßMrjrFHJXr�xX�F<�A`K�P�x����ȯ����T,_��Xm�N
Z�Dr�o릱����cݘk�%��E ��:�fek���N\$ ��ҋ{+2^(kݘڨ����	j&�\_t�vJ�Q�@ģ�v�z	Q�$�
�}�Oj*C@�pC�`Ț�'�{��k:<��q��&�$����;�����޽�c��S�T.dB�2�`�����o(ZR5�Ӈ��ݮ:�H$���X�y����j�T��wj
����.徙}���kTAY��TU8����WKKK�� ֗�|9.��t�ZR�e���D j䥁�2ѩ���8�{��p��I��kv� g{�`�l�%H� ���NfjѠq�:�s��]�{m����p�3�����N;��*�%�����1��;[4zT\fJ&��re<����^܍�CB�5t?����.]r���BI8H�i�4�P�W�(�|�3�`���N]��� !�v����q��<
�?����QX��k�G)�M����ԖO���c�K�k������I.FU��=�YG_��kD���k��n�����
�ljh��&dHۛ�#
��֎m�rA�Am�`~�a`&/�$����bs�����0��˥��6��l�!�1V�� Oͱ̥��#e�����\w��A�1��҈�ҋ�|�����K���_'�E��sCﷀBQ}�\�����I�?k�&/�v��Bv�M��2[R���~mo����z���sf˨L+4ӎ�
�k1�J�hٺ�=]�!�
�Y�����N�ꦢ���0���6�BG�)ׄ6��Kq�& :s��U�#zĝ�țnD��k���{$���}���y:�>,&fn���$b�3�F�T�f6?�������N8^ָ�$B�5(�d��c��g�C�����߂�V��
3'���g�U���O^gm5���@��x��#����_��Pƿ�u`���_	���������Qua�G�0��x�������	� ��)0������{ī�o)9��n]@ݮ�������ӸX21Pm��
H8V:���a��|�ۀSl�)�a��`�
3%�S���'^+�4nq��
W�T%@�m�;7�$#͗`��N`fa1w�C��3�/���%�����P)�झ���	[�]^ܾ���ۋF����ə���t������@����)߿Mw�(g�f{���z��1�~|�H��?�鬈���@���V�܎p�}�?4�3je���^�^��y��pKl%���HΝD��ô�(������myl��2�Uf�sޠSS�Tn#ޜ���>��w%��T���aq�0�P�kk���s�څ[	�91?k�]��Y^��nV��s���Vtm���js{����8�yF����ů�˃������X�����X��E�#f4�Yp���r���\�|��&��/ �S��Ry�~`�R�q���tJVVV&��O��0Ǭ״HGGk����0%�#��VRr�=����$8�mĉ,aW����)�y������W./�/ȁo�`Q�f��,��`&32�	go"�?p�y��V�L`ַ� _8L�rCP��C����U���V�N0����C��D����w��(o�.�l�"rL{[���B��NI�J���"�q�S]�s��G��=�(�yi��7a���B�N�6d�ks�����a����;��C��oa�\<���O��s�7n9!��qV�����P]X:R�)v�����
jY��?˱�@�Mxq]��mp�J� ��L���f�2p7�1\�ূY����tY�OX�@/{
uKEJ��^itgo�v��X����3� ��""t�N9���.���A�~O�p:ل8���(�e| ��h<9�"8��B��M`������CuP~�_���/�����N�֟�V~�}(�KuS����)M�Ť���Ϡo��@�Qx��7�"Vux
j�Cq��uW��x^'�k��l��u���k�l�?��������S L[z�@��;!�]J��)��"E'w�����0x�]��kCE��r�vAX盛�o�?��O P��5���D�p��	a�O�0�9B�� �T��iM�|���[��Wl��5�ƌӉo�D�@���)�խ�	Mt����9�u�E���yi��Ņ��V'>=0���#��!�T�5sZr���������mE���C\���w^�K��x'l%w�t�SS�u�Xf`�~��1E\f���si6�N�G�>jTNT�6��ۧ�po��jGGGb����Adsj"�$z:��{�B��r��>���a<�e�$����p���x��s5����!�9���0m�5�.2�%�z�� Z���Pu��})J��̙x����˰:���W��᥽~ry�_�aY��zJ�"�;dj�i�g��Lk����Tï��A��&۟V�k��=��mi�	�N���;�w�Z��J�sv��ّj�>~�����Y#���{���|j�>�������a�UNv�������q���+�ԸO^���>{�uC�#	�@����N�n���<L��V������e�,����ss�P(�va��֜��'�H�/ Y,����E�/��+�^�v�C�<�mꉹ@2���+]�"��~�KP�5hs�,�/ZlUev�=�����i+�^%�G��}���pa/���Ga�	H��d7S���^�0���d�졉U�v^Vq�`m叫A骏�Щ����(��9g��ʾLf*���R��TH��I$�(��2[��G��:E;�+E��X�O����ɰg,,�����#D��{K��;��B��,�Y4� ����ҴO���R�Tr��a`A��Z	�Kg'\z�^�4�;�,ςb�n��VB5�Q��f�'�0��������^�ϊ��	½��˲r��i*�Z*�s�;
�������U�X��:N�����J.�	�Jm�ވ��E���cK�78�Uw���s*T�*/4B� �_����?`%�׮,���P��o�\���}���G�`~��2} V.�;֠7��~t/��p��f�"�����;v�\~�ͯ���#ĉ�\��;�\~㑮,V�p<b�6ݏU�
v�:��\̮��Y��u�#���Lv�	t�?�</�8lM��aZ,�9��1j,�l�MƁ��cՒS��U`9�H6���|(IP���;*�5��%$��䍃���.���Jl���0`���E����e���!$&8�z^���	O!Z��C:t�=z�(����Ϙ�8�"�`p�����ea+K#�������כ���T&�T�[���L&�771uRyn����+���	����l�p�n�j@#:7�w.�ڝ�K��-����S��4!J�aKH��������?f�1����cR�J�tz�,|�+��lq �l(�W��[�W*NwLaThkiYTayv��d�e_l|���,�ͯ^��ޢ�@�ZW�H7r'K��t7&�/��.}�؍#T��@P�,�С'�Ń6������R�g�d�����u�}������5���.���m�Ɲ�qb^Z
�{0���B��}E!��]�����'��)#�ʷ�^��a�6d��ϗtvuE����<�q�����U�1#��
[���R�u�]��
A:����sNPpp�]Ҍ�0�w�lMq7h%�)J|������w�ޥco*7@7��ߛbq�f�kXCԱ^J��֨Z�o3!�d�)P},,�ſ����x�yԯ�3ն�]˹����]Hk>1��y���9V�8h������a��L�̨�Y����8l�	��Y��oD�K*��P���}���)֟ڮ9�ȘNB���(�N�^i�����7CL����J��$��맢^�4ɟ�Aʤ�*�?���@o�E��/�͊˞<yR��+�ӿ��~G\���������_cƿ�����j��CR��_�`'�k��G�w�<�W*�Y�
���﫽�]��@��?�n��n�0�4�C����Za�e̪��8{�W`� ���/���(ͩ/n��P�b�[�}��k�|-��C��e�c��6H�!�,��Ĳ�^墢H��X(M�%�����MΈGFFV奕�;���=���X�IX��a���6d���;��w#��1[�V��<k+��M�',��{	�v����?�p��U )�@Juφ�:6�
z���huê��| �*(0pޝ�[��{/�ĿW�p3a�N����0�fjj��p�5J���vg�z����k US�Τ�rI�:���ψ*���D���j���+�1�d@\��=��Z�=v]�b+�}�?�k�H+3[_��`(t��ѹC(�ϼ�X������ٻ�{��L�r>�ty5�c�:��������Pيtc��TT�"(
̖�|�;5�֍��"ƹ�艫�*�ހ�u~|�}zL���7q�g\mgF��ޱ�@�3,R'j��Y`� ��,Gk�-o:oi��m�re������-?�����o�D6�]��tn��/����t��i�b�#,��`��B~�X����4�)J���[�e]��|�f[�4������F�@~�B�ʍB�cV���~�Nw�+B�zwd�!R��0����_�f����/������k#Bd�6�i��#��v��x[Ľ��}����M&��ߢ/&\�!0\�u��
o0s�Ql�� SѴ�26CJ��J-�(�p��wnH�^��[	gg~)ĀN���Q��?o��b�|�v�e��n0����k|E�����o8��י��h�; W-?�kY�]�3���v��|�����N���p/A�%O�0���^�Yi���5T�_�4�W� sY![U�xO����9Ō/�>Ü9@��7Њ9���2`��v� �����E��y�o�7H����?�d���[��`�G��������: ��1xZ�;)I������b8W5�dW����L�#���TE������<iψIg��w�Z�R� ��>?2���!O�o���3��d����+�
�T��� �YX� �k5��Y����eh�%8��e�L��^�8U�[����RΗ඗;�F�,�DK=�K�����SӇu{�(�W=;���;7p�f(��ynk�_��<�����9�+���flHI5��.4�)J�6�4da����u�rww�K��,//�
���]q��U�dQ���Nv�q4c뀱�Э��"��7���w7�S���C��A�f������8���#9̒@�`�mh 魗��-t���E�=�ܜb�7����)���=�'�'��&�_~%t(�����l|4�5�;mm����K��p�E��_eÝs0�:�Ւ��Y�r�䮝�j��������Ty��͗��K�ށ���Sg\i�O��G�s"�E��Xa��Z�e8�u3�n��@G�^�I N����*>��蚷�1Q�FLݝ��%CVs���'&e6����oT���cSb勳� Mg��6y8/�Uf�,���J,K��ݨ�jY�z�%E�Ӟ��;�%A7dv3MfUG�ni*#�
CԚϏڀ�x���b�����	���p��]����m��_�pt�&�j�L'c:9RND�I�L`l;��Ҷ�e���Z%9S8/�?��j��}�Z�H@Yg�*�G�<��?ȗ���b7����-�O.3��JB"b�U�~Sj�����<s�ڸҍ�6]�Rŵ�ɾ{�l�>w_¥��x����P}a�4��WZ�3��TB5$AF��W>�3��l�ݱwi�&~<Z ���EW.'�o;����4��g��d��j�p�����HV"[fff���/�aG�-��ɩ�ʉ�#�Sf�5���O��r-�{���t:T�.]X��R�b���?��΋�nooW���5�̜ P�τ�lT=������~E���*��1�`�ҟP�^7������g�����\�!-�{�o�ӷ�5O��8JZ��e>Zo�Ӫ�ԃ6����te9��B��tj*�B`zr��c�0>��}�ǻ��sL:?8�����u/������d	Ď�z�X�;�������^g>����춾Ɯx�����\5\�)c��7� ��������G�U`�
-��zVR�Oh+).��M�@.L�#�MLLT���*���"@o?@�ܻ�����V�����ϧ2�E��H�I��;��G}D����C�Њ����o�g�y�&�*I�*,rZ�	sI�ύt`�>��Ϟm��[o8YE! �SR	�*�׃��/y� v�2�`[�ƚ��$��(p�7?\�ɾ`���3-֝6y]��Zځ\c�8/������F�zJ��c0�N�,�{�z��2�Q�0�q���Tؓ�G:����Oܜ��k�8�@K����h/��bL�ē�[�me�0��}RJ`���-���sQѹ�Oݺ{*T�t^t5�T|zJRj��ʉ,sb?��T׽_綍(ܛ�j���L�kH���T*;�6S�l���#��[b$ ��I)0��ውR�?9(Kw�
B��T>�L���?�S v���k��I�TlbjF8P�4��v��14�����[v���+��k���8��R����P��_���h4�#i�9���IW�&�N�Ɗ"▛�"�<��HO.M�k�ԉG��I���=,�TD���n�Y�G&~��;񂗳��j�-~s��?���7�'���7��8�Y7P��h�,�K6�%�%��D�C��O`��L!��6��d���V��8����B��8��򪢰�b�i�i�L&N�u�$�a62#�`��N�i���7�G���]� ���؇\&0����_�ϱ�^������������}5kzΙ_g��� ���Wق�}U��f�.܋�p"�w��y��P�~ۦ�g}_g��n�����&�m���~��>L DK3�� m>0!��Gw�%�_sV3��u�P�l�ٟ��ͷ�x�,v�GV:�{"'櫞�T7Z���D���^T�'�Ɨ�V>�,�/��2AD���¬2�{�rPf��e���bn�j���F9Gic!�ɓ��o�ic��,g/KD��E��@�q��� �8ƾ�g�\-�Me��TV(���v�Ut�Cj�c�Q�H��O���'�V�*3#���+��W�:��Y������jX:�[��p}��e����\+L��vL�ǡ���-[c����@A��2؍0@$R{�">AҲ�Z��r�e���"��/b@���`���q3��骹@�e��w��2�����l���.�y2��S������A�,�m��ڗ�S���'e��Axl��C{��kim���~�ʪ帞���3C,v��S ���0��!I����:�����P� ���%1�n�͕D<�-�SZ�"߫f�����GQ[l+p�)|��~O�.���O:��i?�H��fP+���O~���2น�����+��[[#��2��F���'vgpJ�N��"���<|D��Y��(��5W|�6AC���!tSu�5|�+'<�����6H���tϨ������Y��?��:8�d���={e���� ����]H�W曈�! c�J~�mՌ�ԕ]l>�߸�#�	.��]!$��wǂ�"������@�iY��j��c]e�!�<<�u8~��~x�"Z
d�C�,�l��J�6T w��WrҜ �U.W�E�����:�x%E-���z��{��S��G�3�hN|:�g��Tk�:�)�♿w���Z��f	�$�S�N�qhW�v�Ŧ�͡��o��mx�.!Q���������8�
������{���w�Oj��'���T�9�B�����E�:��/�{g�i}�g�/��?m|�	�əŶ�����Gc5��˟7��k��=s��6�.���w�lK���V���C�(H���K~i2�������V�ϯ��zy�'o�jw���<�P�TP"[���u �;8�Z;�::T�G�[~Wyv����9�ف_�p	т�;����W�H��p%�G����Q���EPAZ��o�j�*�B�x��Iw*�z;%X���a���M�b^j ���S�E8��L�d��%ĊD�����sX���k𻀄��1<d�'��=3�A�#�z����j>k��{$)Fh+X3�_Ce��]��AM@z���<B�xKI�Xx�#"Kc��pޠ="���CWr7^f�r�&�\ ��;�z�IX�D�ajn�t��(��E��#z=�����w��Q���KX
���o)n���4˦����ꭻ��y��JV<E4ō���9l�-����TVN����>j�hH���{���A���Q�Ұ�Z�!��Ȑbj\v�ۚD�r�=���.3ŕ>~��Ȇ����+�}���bhc��(�7��Nu����F��yP����%��,��ІDE������D���L���P�U`�6Mc�UW�oZ��̢B/��i3�qX./Mx�Υ�ƶḌ���ڦɝ_T����i���g���$\�_��h|aڧ)�?�g��95��M�8�T����>B�Cj a�;~�)���}�Z��d���Q#�i�FmX�jZ�#@�����츖��R_Pz/�P�T@~�H�Ix�a�?��X$�Kj�Mg���ڵk�:15<a a9a t���w�QՉ�Sjg̏Tn =��֞vmM#�_�����_��`/aLL�\8���Ӄ`��@���9�Ņ����Ye�mO�l*�]x�'oQ��<��-4�ľ��ե���)7@#��/v��⒒z���h<����������k^Y��bM�5=VcE�&�֒o��"��N�`��?���H������m��2C|�n���Ë�\���̳iP��~-/�w9纕��<�f�.��OdP e�=�7���~��KSD[���1×�\c�r��f�;5�Q�V E���w�b�j%/�Q��/?}�O6p��_Ɇ4�gʑM����ƛ��,�ih�^�u���/�T�qP�=�fց�丸����:G~�Ƥ)/�%��e�4TϏKu^!�ѼKW-���<���2m��ψwL�)�������,�����=�V�$�E��΃�m;��Dw53���ܝa�CA��������wj����ȇ���	]QZO �������3#_�N��w��7�a�z]����	�ࠠ��ϟ?����	��)��j���$��U-��AmJ|���m�G��,�p�#kr�����ˁ%ʝ���lA�+$;ʡJ�*�����ǟQ1O�Y��L�؍�5�9^>"�H����0�\t讃miǿ}V��g	!l%-���5-��[@v�������*���g)���,1�(��i�d =�(�{v���DJ,��A��׹���Px�gڨԏ���{�[����h�]�俈��~c�ɩ����="ԟrb�%���QH�����V�z ��c&g���FFF}!@Ӵ�],�w�"�]R�y�L�a�;�p�'�Hq�����Ι��k�����&挱z�S��� n3 0�G�	�0Y��6�DćPb�O˼��N��ߖ��u��	"|����s��O?�	r���<=>~	S
�C� �� �XA��"q�B-�HR��΀��چ���
���}%wOE�ӟ�L�j?�1��[4;��2P�kl�ŀ�HP��G�̙`�DSvPÂ�h�Tא�=�I	Xnj��{y|D�'yflW�8Zs��R�.HA�|�yN+(e6��h*���(��d]c��]j������� �'���S}e5CB��S�� g��eM�w��A�i	cM�_���3wB�5����:D����Y뫕[�KJl/qo_f�[lK��̜�An�|�in�(�Q~�c��f9m������O�+�G�Z	o"c��"�[�tPkY�L�U}f�4	,���:˒�Yb�OXp�<$k���2�;}Q�>@�PjR���}[��~^r��Y~�΃�Nv)��'���~��{���u�3���8�0�h�2�oÚ<2_zؤ�Oi�����SuV޺;��5�;����3��e�+�>�5��3�.:Z�t��%���Dqgg���Ҏ��j9���,~�^ ZDI%�37�|�_��|L ]s��Q}$�}I��U�O�7)�݈��p3�����A�wD$T����`���T*綽gFvF��|�DFKK�Bb툟 �KmA���`�,>+̓�/ׁc-���C��^��w����?M�^���0�Ը!��[P��[����ڹ;�S�yi�I�8��;��� [��CPF�u[��������aP.-S}���4fnz�5��K��]��s�������f���ڐX��u�/Fk�@qBz
�]�`lV�n�m�:�[f(��ù�����\���]0��~^�37"
�@���ן�΀U2�⮫u%@�^ P���'1hEl��o�%�$�6T��YBQ{*�Ea�Y�������{ a���npj�	��넷�/5��)�[�z�$J�}�lQ��L!�}���ߨu��J63ǢZ��g6{�^�i���~'��N�:�]����'���o�U`�{���l�����qcO�>�݀.�e/N}�+�¹B@���6�?J�T7��y�* ��\hY
�Ö~�E�#��1L,������2*� 2�d������@�07Hf-KҜ��Bم��f�T��^�� ��|���i�����l\dkɭ��p�'�Z%@�m"��|�`�?������h@\PAr�@kX'�򧥋��*LrZ��If���8���J��L.���I�S��Y7����#:?�:�ɬ[�4�&/	^9j��S�8�L�`�A<���eI�� T��C��ޔ�����<�}]ϼ�ނ��m+ùw�7��S�X���a�(���b�[a�N���h������i��H��"�� �ςh��
�a��������5�@,Ő��ݥ����Rw#ŏ�1cu�|%��ږ��'|��H>���л`�X������MP��5~ĝ�q���[A�*��	8�6xA:5���������u�����o�:{�K�ڊ�m7�\j�]��!�]%���P2��Kr�M��"�M�vkQ4(M���&]�&+CaL��eH	�眷�����k��s��<���������Ґ��K��M�$��Aw���i{b����`��@-���q$�kq�e!�b���6��4���t�������_�ΗFVg"6S�װ~Ov�hY��?�a/@�|���LFM!$³�#��˿#����332���o� $ j�L�{�!�z��"S3H�T�K_.L�
�vg��;V�Ul�{�\Cgv��!�z$��Xŷ���⮐�v�+V�&�v���u��V�V�N�{r~� �x
hPKR4cC���Ɉz
������Q'�G��J_+4A�\V�e�ҹ��D;w������OY����@jF�~aKw���
�X�R?/T�XH3�5���L$�#�(R�=�.q�?
P�_�&�2�a]Q��(RH�03�~V�{��6����� 矠����I��|�X��Xо��d&/��lc���ެ'LG�%��z�y�����W[�S�rj�{F|�o�W7|��jii�-�;��G�9�@Y^R��yx���Cg�f�#��:O3��kb��H�m�`Ψ����u�1��9���(��npKV�+c`��I�*�\.ٓ'���[����S��D���H��#`:=6?ڕ��d���.6����H�$�4<�m���7�t�,��W-7�����TA�7��i%e���[�6Az�J�V�t|F�	-:��R0�$�(�&S�*�B5p�5��[x� %��|�C�K���z%s�
��0{RZW���Y���k�S��@�y�͠��!�'�%�b���}�m׸���߂k��sZ	�
�~�ȓR���G�TQ�x�/n��,YJ����;�DZ�h}}����:�t�U��ji��_��%xÆ�����hZ�B�mj�]�h�U��r�^䠘��2z��|����Ѫ�����j�d_�n����WK�}�����'a*��E	��9���VVU���}�#(nK��"5�`Ah�U��o���1/�������"�I��}�T��8A�%�ۨ���|e���%��oq6��|l%��+ӆ��ž|�޺�њ'L�F��7���S��[X)GӤ��ܲ;��:���m�L�t?b"l����7MWԉu�0��}���gtRx��ѵ=+Ge���po
Z�D }w5���q����� [:����?��#t�755��:U��->���t���1���dYXm�D����|�� ֢��nk4�@�8��Ldk���N���V��N�����:��H��=NdU
{�A� �Lu�|ŋ��������>�>��Q��.1����;�z�Dښځ��+����+#��y�5��<0߰�H�ڹ�xT���ka�ͧ=�rU-C�1��.���]Ƙ����#��sd� ����<JC)���v��5��c,�f������S�tDai���?dS+��-�'����ԉ�R��r�e�"4*�����G7�� st�o�#4�揦��U�]�wS���(�ܻ� VTGQ�ea��OeБ��?���`�Q��8Zc3�{\��1p�_�U�)�	Y�*���:F��}��)���IB��Y�����ƶ�����@*�Q��W���Z�T�_�xa:���g�)���mu+�%��@�;A�c�͆�;xo���b���c|��96
�(m
la��2ާ���)�@�S�������Ĝ�5-�ãr;�ܟ?8��2����^a@�ru~s��0;���ի��H��L�	�'@����&�FcZ*�詶	].���,Sr�:k�>���s�S�`z';�Wbb":�YA� 2�����ʗ(qgqF�́E�h�N69�ri��P93���[�/��BW�@L:�Zj_�^E��o�X�ʅ���V#�Ɠ�y�+E�A�Z��c��^o�=߰��XA`vbD=��%0�:%�S_���gl�]� \W�ŕ��J]�ڶlҦv���u��C���ZrBT��=w�0����۫]�\H����#,���GO.(1�����C�	iM1�jM���9��9�w_\���a0��Ӗ��Hti�.v4�b������#b�I����>wa�貈��w����[Fi��OO:�wQ(-�����.�*�p[�fϘ�?B�4-�]�-#��a��s^��dGVEch�>�
(���W@�q�L���]!a;x�P捊3Q���x��&sK-�Xl>g>5���p[�ߪ�Ӡ���ʋN���TQַ�0�3\�o^6�Y��YI�#DQQ�#A�ԁ�(3�zmkFq1`,i	 ���%9�F~q[��Őa�����Y �� �y��ǧ�b@Υ�;ܣ������Z�����7�0H��iK�OP�Z�	2Qr�in��~(�w��k���K�09re��f���.9�$d���H��ɱ�'Ն~w�y�V��.H'�Y	�G!�wzݗ?��5���������T��/%W�S��TPi6��'�T'���F��݅���#�	�_Q�ָ�xi��Ps�W��h@�)�{h�whm���zuJ���ܬ�0�]^c��9�o��]?��i�~� %3 ����v�2��I>Ƹgl鷪��g��(VL�Ku�_��Ϯ�M��T�zFa�
Q��hP ����ɗ��g3���mlfڰ��W3�!����c�gT��H���Ooo�x��AȾc���b-��7.H+O.v,���N��㪻h0�ka�Ç�>�����y�FUP���u���В;�!�N�.�
�T:���	����8�u@E��db�¸XWGgj@��N�U����;)e:�u�8��oe�wW,;u���Ө1���
�)��0���7���%�";J��,�,�6���
�x�A&C1�n�I/�0?�mGt�:d�a���V酉���]�[M��Y���y�>�)c����s?��F�+��V49��a���w$V�j�Z���5\�jv�Ü��
i���hٟ��i����<��^�����s���J��]�l����tE���{��)�eG��i����1��`��I��(��Wv���>��Z�v
�HA�Œ�hS��Aȧ���4`e���;_��_Z3S�C�d�Ξ��m������0�.�����#�f(|{M ��T�Z�Q��{�/uȌ��I�!uy)쀬�B�|G^�9�E�r��!�!����N�� =�v��=� k=��f1 ~�*��5ioksKv��GH������|N^ԙ�Ǌ�`X�� Ai�O]d2~t���4$8�%ga��v��i�R	J-�+���q�s���"���u�u2��C��Q~�GC��5J ^�tF�3�W�VF{P
�3.:%�=_p�g�bj�6r�ܬ$�pN��F��B}r�>)��?L�n�Q� ��p|"=�2���E� ��Q6�	ɳ��M��|��o!�*���Ѥk��9���qJ�iK�!����ʼJ�	e�癛��u�$�P<��������
jg�Ƀm�q�hcƨ-�tHS�l�?��5$��\ȱZ����gؼp�"�oԓ�_����(���j-[��°'Q�[h⭡�u���@�҅(�/�̤��$�ѐ�8��j�������Hh�Ը��%��:c�Y��|p]ѳ"4��t�/9�Ȳ�L~U�`l?�§M=ى���=.�nɊ�x�~~S�A�)��	)�L��3���^�i_�ZO��wl����!%�n��=��x��fy쾵K=6�C�J�C���_2�h��p�Tx@.(���G�V�{���9}�m=�!���7vAN��	�"]�4���C/�-��VF-v�]���o���YD����|ބ_P��]��/}�=#���9�:�� Z�h	*�ĕ\�$�Y�zH ��։/8=�H�a#2쾆HV'����u�胶g]���̍�xI�!z��Kڻ�uB�q���h|>��"���<2T����a>-��.�?��=��S��T^�ۇ����]j�w���ť�(�Ԯ�3sD��S�>�x�F�.��h{g��f^r@!\^vgp�'�0U^��și1���j���nI�*�߮�1�к:G�'�3��cB��N\i�`
ŭ=����P��!���pg[ ���N�@�\.��h9DGSn�M,%����D\;�
'&r�/�x���L���^ȕ#��^ˈ�O�kz���\�d�P�_�pT)^[�
Uz��'�D!����Ј����9ROV��ݢ���~��{ٟ��آ*p�xϩ ��c
3�/�4�A*��wAk4�W,=�����<�!��`2J*��!�@�b�
�Ə?/e3�! ��Ͷn3���[WS�<!>�0E�2#�!-XH��~tD�
���mޢ��f��O�v�l��<�d�i#�jM�	e�X�rL�#�X ih-q�;C��6��m9
�S���״T�y�:���βu��%��W�c�����`F"˸���c4z&:vƧ��m/�\������i�Q��o?s�_Q�P���V�9g����eG��/���r���{/揭��w�Y�l�9NM2g��ymǘ�[c#�ё7�oDG�X]�H�"��s�Y�	���T���Dev�q��Ϛ�Ɣ�
2���I H�����X]�`��rp9��?�)[���"u�R������v��R�_�"M K6&|�{]�Q�Ԁ�iP���d3�����
Ъ���G�:ѲL��i���v΀���c\�8@�@�������S흒�-���M��}�h�@�P��Lsǉ��@�Ƨ/�l�M���	�hj�ܹ���:vfW��{A���c���'��T�Q6��*��@x��������=��>Q)jDc9Ʒ�[-���x�c�S\�k]T��>���$.��(Z�q���s4-Ɔ���Y�r���x B�%r��!�S:�?k�
��-0�c�O�&����� ���O����&Hy%.��,:m��J�xCW���x�០}in8ȃ��	��@�$@�՛���[�����:&���;D�?�n��P�� �k{0 �|;Ϭ�q٧�0.0���='��?�w\O~��;�@d��6�Rd���!���lH!�m��9n�Ĕ�%_�qH$2�ᇆ�<�L����m����G�\�(�9m.�Ml<rRMt�˽��{����8�Kjg�4�vB�µ��9��Z��g��w�ƕ-G��)�v�A]WQ<�6R#8B��]=u̓�G@����e=C7�/3� �ė�s����
��9!;�K73sQ�h���f��s���8K�Z��ݻw�8T 7_�6	�ѐAâ���w�!{5��z�	�n��2Ch��.`�0DY�ה����HS�j�-`���8�ܲI ����������xT�J��54,���[���HcI�Sr�A�+_���-�	iXK�ڠ�a?�گͩx�8����m�u�k�g֎���c�w�d�-g�e�w+�	ly������
׼ ��A���A�"IJ��;��>QU��2q��qS���J�u�@�|��D^�F0��f��HuJ����>s���9'Ba~zq�������"�3�b�e;x&!%lk���\��ۏ���YZ'�����7 `��(����w�wG���6�]�#4y����-���_УV�U���p+L��@D�1��d��tWs"���JU�.�l�����h���ϟ:}����-8ܒ:g'�����$ݜ8�興w8S	CW�f�FL�r7z�&����晗OX�sb�o_�ۮRy���� �	�pEEeeT/iMtS�+�q�����c|}�sU��m�����(H�\�[��M�]d�5����b�5�]����+Z.w<�S�M�2�(�*N�1�����h��P'��������M��ȑD��E{
m(�#�o���i^'狎��ks|��h��|hrmC{���o�������I����nx	���ݹ�v%��ճj��{��o���&����3K��x�R��0/��qe:��v�PD��A�|8��{�ft3���lr�щ��!n��J�w)}}}J�nJ��}�R�9��#�@�{p�]n��T��5ϛMB*~�M�|��ZY���u/��߲�_�Z�^sIh��JeC���o� v �pM���5�
�c����z'��~ym�׋�+�@@��/CG�b³U�%b7w0���C���\�)Е�|��&��k�e�*�m-xx�]ځ����3�n����t� �u��K�*����� �}��o� �¾��\Y�yK|	�z+��z����r���=8��j��N m]c����R��V���d���'p�s	2���6��H��9_����Ge%�&1��k����P*T´G ����vn��n�9��;���?@�Z��ܪ���T�Ӯɣ�d�(`9O�J�X��W��9�rǪN=r���Y70�5�+Zx�O/mN[���#��.����8�v��}ϵ)ٷVf�Ǡ�s}�H��f��F��a�@�Id��Ӡ�����G����C���D�U���Є�B�D@!��QX.}�Б�¶Z�m~PK�W���B����d����'�0`��T��w��\"�������&�y#�i2�������c�*�Y8*s�V��㕿�jRl̳$�����D��S�SU�Gk��)�.�ۄJ���`�9����zA��G8��� �G&�$b��9�w#�r�׏ʚI���9zB���:Z��2��~L`�(�D�>�Ԫ��_/K#@^i�"�#��
�&��6��{�	*���H=��I��R�kbЍ�y�)�84򏟻m�⅄�ap꪿�,"�/��M�-��
��O��� �*H���0 J��:�7@�"rr����7�/pOv:�
m`&�&�c�pa�I��mG��x���ԉ�p���
���5_֮��t��9�� I��6��7o>�@p�NM���`�zd<�߶@�T{\Z���XHP�%��u�7�]�9ҟWƝ��Z_�,y�ie�\]�}���m!zPe=�/������m�W�����t�-:a�G^���0{;�5��W��1˂^tޟq_���wlA��{#�F[V�ҹ-N)dGF*Ȩ(L���}^�	�����3���W`bj@+6�^��,�xx�S�x�;��l�:�v�L��@�Z�dǧg�>�T��_�í�tw��?3�GD�*�,p^|\U~^ }��h5���	z�PR����ɳ��d�+�.	3��{��A$�-t)�_;H ��h)����*������ԍ�?G���;hai�0��*O�L��\n�0v��۷�x� ��˹rg�s��/�ޭ��+��A���)����`�t%H�怪�o�oF���G�Ңg�$%%UӨ������U��x�%;�P�}ݱ��'��9�y7�6D�n@U�A��>(��uߤ�/
S�WF2|��?}���l�����Հ�7K72��(��w��Bt�/���8�a�ϴ�W<��Q����n��� ٢�S� z�%�ː*
�������?����6���\r�V5u��A!��� :��PR����G��X)k���tM=�I�$'�c�yИ��]�KB��|�]��5B��m�m��*���5�b�m�|��Æ��+ڍG,h��M���r�O��RY�Zh�M�@��,��G����~'��a�F��Ի������
GB�jEq�#��*-�T��Wo�l�2c)��ro��g��|ǚ����W$�����J��9Bc�E��ָ �X�X�x�Ω����TV�~hM��MN����'�B<�Ğ���I�%��"�d���|A�C{kO@,�T�3PYJ�ڷ'/`0�	�w��M��-�׿#��Pt9i"w|g�����}��H/b�g�i��]E��!��z�W��Ya9�5�{�e�.vqaT��`ٳީ�b��y	�y3���;8�C[�}̩���@�[�vP�]*�)Rf�a���RnM7c�����k`�Gt����e��h�L4�["�z��'��n�; [UlE��q:{AL����>�B彶���Lmk|��ym�ď迊�7���������e�!��=`?1֠�� m��$;��BZ�h�g7�����ĭ�EAe�n���+���
&�y��իj|��(	��b�5��B{�g^�i�n�(���smD�qvno|����KC*�M�gcc�6~�4��I}ڌ���KlP&d�1C��
��;�/����4�-�U�t�t�Kp��:�%��zs�b"�w�`6����_P'}v�w��ڠ=#j(�)N�&�S8�����*�C;���r�پI℣i��'��h��:��.��i��˞�Z�3+����>��==
�R�F��O}���E��ND�*Zڠ}5��-�ͧ@s<�%�U�E&{ OBHѽc|MJ�I�i��m|:=C�<8v^��P2���m�o��n�mv��&�<����,Օ��סʃH�!R���~+F��{�^�Յ�i��
�D2S��N�A�7���xx��;�m^��'��d't�BєqPS��:�3 �s$���1^�j<�Q�	3����E��+�D�bҩ��Ԧ��\;}����M ��'��?���v5U{^�W�`pd��/�ŏ��n4YgŢX�xV��%��h��채2sy��g�>���7�N�S��=�ro_��k��4�v9yO�uvr
������9o�:#3�*IM����9�]�C���C~rwt9�d�'�钠��Y�K7�_f)L~����ۤ���w�Bͮ9Ƕ��Q��	z��c�OU\�yU}{,K��5C�v�������i��ڑW�%;gƮ�H_�q�Gqh5��ؓ��p1'u�C�~�^MLT��!�+?T,o��?v�����5���C�e4�e��=3#?��=��6Xix6/[;g�WH�$R&ZSߏN�D��+^��;�3���u���e�'���`&�m���oB5Qh�D�jr[�����'��W\���&��h��m�5�wzx�c�^��F~MӘqzk�z�9�,~ґg���G�9|_c�[Ԡ��+D+O�D~��[6+�qS��M��FJ��X�؍�C�YrK�#T�UL�
�M�u��΁��hC�Nۈ�����3�@H�������wɜ�,�[���a��M�b<�܀�H��p��o������({�+��B������mbpk}���!��$�GE�2Ԉ�,~��k�E�Sd��W###6x{UQbf~~>��u~1/U#��0 ������r��o2!X
!R�z���	���j��?��C8���*��0s�M]4�;�/�BU�2��ߠ���)e���S�y<���Dj��L�g�Q9�ӟQ��vi�q�*O{W�>�`*r���q�I���u6�Zę*��u��z�ם9/9�4�l�E+�)/<i�{&6����������(g�����-�6� T�5=8j��D ]����{i���f��Gb[�����c��I��	��SOC46�D�i,4*j�Z���^�������Hk��L(��"��ڔ^�	�ƺ;���m�M��������R�q8ףm��N0Ζ����@�L���\�xAV�j��*>�r���/SX	Uo�8�$\��@f�q�oB�t1�K�s":z�J��}�R/K�{�RU6쐈/.iS!�?U��pD�T��XV׻����F�(�R��O�|{�r�����n,i__��jT
_�}�hZ�A�&�Pg3��V�
!x���ՉCFRw����<}��̖\�1�����8�/f���<���)�D.�X�R!2�aɭ-@ޫ�nd�����JT$1t�^�l]�]$�C�
Z�LN`wB;��2;Y�޺� }�P���d��j}$ґs@�{fW��T�N{��S	��� �S_��+i�js�!�M����*��m���޳��dj6$�np�;=,�<���}7�@W9�vĩJ�罄�1�{���7���&x�yԘ�7*꽺�?�4~��W���B��$���7o�,����@��|��[��c�g��~�~CK�v��l�w�j(G�$LWzvr#���)���E��x�MH��n��zC�4���G�iي^ǂd��O��d7�j��"�e���h�f��j�B�m��!�K�U��;#�#a'�j�*�0��ȯ��׳��(I�p��mM����lՂ������0_0�t��PZN�8�a%�_�
r���j�8�7�?緜WKpy���S�"�If���i���S�S�ހx6R*�;<��5U�z��tq������h]�)I��9�Ӱ]8�e�e�M��M��eO�^A��>�:�[=+�d<Zop�p�P������SN��.>�M�������*qA]t{�ɹ�$���:�N@د�`���{K��#ϲ�t�s^�F���%}Gu'{�X@'��c�{dV��'h�cd�&Fٳ�%�I������L��gBKZ�����ai؟�}�+;�?��dz_�Y+�j�[H��M`��\�S�U���vѩ�H�c�)��k�A{��h��S�C��z�Z���hf�T	␭�`u�$�D��ˡ�m�hL����-�����W���[kP^��(�����=�����v{�/Q�����yhM[ܭ2�S�zw�y^x{��vT���ÞR^�TG�3�'}w�a1��>: �N�f��s8S3���NɵlAG�(�f�C���HxZ�2R��ц�����;:H߭�E_9�{X��H���Po�GE.�����#(�"�^���ŶO�z��/��9���u�.�Y��yV0��bj5m�4y�n��&9�����;WT囷�D�7��B1�����s���k�Ӕ�"Ϥ��uʋNU��k� ��1����;3���D<�`:�[�7K������C�E������	��6���W���;j"�1��Jp��
�UT��!4)|��?����_��D��D��ֲ�7�fe>oL�Voϓ����GiJ�=nCv��y��ф���Ԩ��W,=;�������EM
�{s����S� RG�{U�{RU����U�V����I؛��w����N�� '��;�x��3�v-�C6�ɕd>#�s�lL�''`.�]����t���w�q��E���Y���b�m#<��֭R��Y�o�l�q<.�]4�o��w��Cќ�������I Kk�ǃ����qܣDZp����n�ᚭ[�ą��m����n�C_塟�ۑdі.��*��dv�6�r��c�j�rt_�z���W�}�2dꡫ�=Ws�Jp�BWd�Ѥ.��3�ɔ[^ ����h��mnX�K� ����D�
W6��es�:�yz��k]n!�� �q�N�<�0�i��8T�ǘ�'r��@1	q�a������3RhFVS���s��׸��n��=�����2�C�(]����mZ��~�c�A#z�vptt�#*���߇��m4�_�QS&誦� ��-�p*�#�˟��K�kh^i9d���r?B8=*6����$9�յ�z ��&�I����Օ��˱#�<�I��O�k
���rձ��;��Ӟ�)�NY����C����K(����ڠ�Gb�ϑq�U��8|0à=�R�,���=�!�Y�M�XtJ(�h�X���h�^�$ONJϥ�c?�����<��O,�є���`[��?�<��� F�vl�&4E��p�y���Э�-2����%��k�L��"�ſ?�-ɜ�&r�?���M8��M�A�n$���7ԧ�:��z[vS;�\Y����׬^
=P@���,�>��L�X&�_�Z��Tu���W�3��}2Õ="7��]jzX�v�	M�(|o�O,
x>��L���aƔ�H���
�ė�\�;��W9���O�]��Cl�=�5�� ����}l:�+]]]	~� WW�%�3\�AS�"B����݆x4��=�#��0������%}�G4�����C��
���&'������o�OԱ���h���r#�U�@>��h�����(�y��� k�^a� ]�ӟ�~��˰����Q�^!�����0@ލ<��o0v��$���4
f�0���d����fM}��8��n,�)�ŧU���� lt��y�3~�頀7��9i�c?�2����Bȴ�7�H�#eO!��"��"IZѠ�2�_�&W���7o���3��x&4���Hcdu���� ��G�߿OV:u��!R�!�bChd�Oi��|��	lL�#?�XuMP�O؂��|>o���=�s~�%x�+'u)�:�$l�o4{xxT�`����{����24�w8���|�K�2�G?;��	8���nN�������^�|AHӿ|���l"jz�K��"��W��@����O�ɜ"����Y{m9�3J��&9~x�"SD�h���1~1��2��4�����U_H=�$��/���/��3j*�3��*7��4�J�.�|/��K��.��7<���z���~RuU����K�v0ޢbִ'i9�rf��g�.����A������m�8�=�(�!y�!���hᎼ��=fs@�*;��.�U��fS��~y(&�<N�I�ܴՓ8�>�f�Rb�%hn!n�A4�wE�&z lEcĸ��w���@��H��`a��W�n��0�C�$	��5�~��C�'�ji�}�v�xIa
)�'ZvgDՁ�&w��B����æv�x ʝ�٢�c��6�O8vN�b�0��A>���|��3�",��mE+�UO}{�J��Ҥ(���{<��@9rR��L)Z��q�L�H\�����*l�_`�V̵K�+m�f�e���h����ÌM��J�GR�w}��\ׁ4��1��W��C1D�pV>���p��=��:���T��(N�5"�D�}��Xxl3�4��ox��j'{��?��ag�����sT�����n7{����k�M0-J9*���l^Z��_��}�˗�'o�%J�Ю(��cSI���
��6�h� ]��{ܗ�&�~|���:��;ft�9Ry���/�5J�E������VM|�$v���S��@1f'BW���T�k�G��͞���K�P�� �Z$B����ۣ^	��uD�sKT��}����t��DS\��t��8�2�W�&�2&|����9�|�:{�Z\O�LLJ�1G�Q�s�\���G��'�j!n�(Q�,�$�<#�y��E�B�RW�DH���>.;L� �p0+x���\-D¹Â���9��b���6u-�#l�Q;q�����G㶚�Ł`�'2jԶ��
��,H�T�9��/\r�dEL~U,�R��Aѡ�7��%r8��u��D�&�-���ы��#� ��t�3�d�%��{��a�Uh�(��8A.7i��v�)xޫ�7@бԈP�lo����8h)E�%�mW�g�+;��th�x�]-J���Uj9{T����P�q����/t����t3����&vj]7y+_�=0�R�s~	h ?�؛܀KQ���G�Ll��|������/�.�{I�@�ܳy��uاȀ؀�6��}�ҵ�����
H�(n���{�����ע&��j\�j����$�~��|}�=�rp!��@OS�p�@���2̅:�e%���%��B�������nD�k�,=]@���}�i=L��-���� �;�����wH�����Fo�t�736�ʱ/��MLG�.�=��r���s�(�߼qꔑWK�l_�f4cn�#�e���k�����h�ɗ�t�w�5%xFxM����j�����&Z!��AX�tA�`˛�1q���^�X9�/��i��U���Ǎi���3�/$�6Z&�<#+k�Ͳ�ծ���=:�6���+h����;>�v�L�!�S����Κ�(wlr�z����E�G���{�ծ�y+;0A���g��><��&	�(���H/��J�F�$#Q�&cպ�Ca���1�:�2}���>��V��o�n�=u��O�6} ���>>>3�����f�,�`���"�B;�;~^�J��M$-~�~w���=�����9��\����Y�}!����8s�%�h����q}����(�6XM�mMie%�n{����r�M�щX^a�(�6L�n0�/}D�!�)���8e�Gn��#	�l�{\%Ϗ�� s}�j?�m$U�t��c�ܩ_ �^�L��y(�p}l���nz�R�iU����HK��ڋ�C9Ż�0��E�q���Τ�%�h}~���Y�:0֊���X5l.F�G� �s���=1	����91�L������44��D{��'T����Z��^���`<JQ�+a�!��Ρ#�L�`���d�]$��&G�<%	��FMM���Ĩ���l D�75���nBkt�:B��'����0�>�;ohhz�'x��d鯩=F�����]g�K5�x�^�ul�ϣi�9�*Љ���W�Z�ć7���nu(fب����W��X�l�����P���}g��.y�\�Җ�C��zn�T��ccc����2�|T;4���C_��'CB�νV��3T*������|�����=f������jK��B��hZ�n�ki�.�ѡ�mgFބ��T���LӦ��)��_��s��r�n�ЀΡ��C멝zy�=��Ao�����lg��N]F�g������R[�[�:�?-/<��{`��i9�R1��A�<������0I���V\�:i�R��T�"F����g�'x��6�g��o������ڗs3#^{  p��+/�h�8>�h��a֞Pb�.Ȫ3Ҟ�X�q��-~�"{;x�L����[F��kuN�^��Z�M8�fה�OB&�������t��z�:_r���_�����3���S����
Y��;M:EK)����S�Mm�^;�~[���.�nE�0T��0��mO���ݘ�b��.��/�%䦣2���w0b��������?�o��H�K�jy%K�Τ�k�'ԳF��`D`��g"��B)3��ee�34����jMiv��W7����h�(�PZN,�ptd2)�(�+�nv���X����=Z�߱v�
pf&8�qP��o#F��$6�Y]�Z��}��}��I[��+��xn)��hC��9e��kߧ��U�0�t_;��f���h9x\�k\��|Q�>}�Pp�f<rF���.BQP�J�\��d���Ka�]-J% ��T��2يk@�\�,2��Q�_������A1��g��D)�*�yC��/�	i�wV�$��4g��p���ݟր뉶 �𧦕ձ�U;!HR�]L	Y���}m������3-�����wO<��n�i��jW՚����}�
���$kDQ��^�J�<J����K[ƣ��z�u2!�w�q*f��߇��KZ��Q�P�	�ড়P1� OF�L�u�NL�}�����Ʋ�5��Q*�~�dz^�f�q�{F�<�3�[����B ��r�C#r5�o�^	�g����!�dx��-��PL݅�>}4�x z|��M~�X�$Z��� D���b3xHZ<^���ŜߝX�LvP0�ۢ�у����|��v�s] >-�P�Nk�5g�­kK�����~�#}X��q�ͮ��>��[�%g3�4=������{���5Ԙ.���
��������Z�:�,�O@��q�'��ح�y��I�:Ѓ�z�.2�l6�����I��[d�-��&� ��j��Z]1��Sy�p�ƕ�;a�[�q�ѤL������<�5��~ק�GM�8mn���_�l&��-����_H /�����L�����k�)ʘ�߫���z�SyWHT���q�C��X&q�}��uk��J��ϕ�~K�A�PL-��lWd^ý]on��8�T.��~d���1�(�(d�S�&Ɋz��c/��W�<틈aQס7� �-F��m	$�͗R��$>���Ӓz�^��K�xe��W�W9��_S��Y�`��3��|���㹖ȖD�� Gt���QV�: ���R�P���=��:��)
}�<����ѡ�o�_k'&&lJ����i<k=�n%�D�6��l�Y5����+���s�BA2:��z��W���Y���*.�utC_f�?��
�~�)��P%�K���pV����=��"'�EVw�x�v��}j� �Gvy�t�o[c���,���Tn�⢀&U��Z]Q�rސBV��W�,���)ˀ!�c��2���01��'�($�I^�����R)A��@*\َ{CE����7 �+�{�7ܕ�(+~>�jG�υ�'<Xum�f+PE�-���^�΄쟸A�p��3Q/��}�������S^��Ρ���ה��k�Z��0�Ïo�Ү��s
_�����*B��Z�4���3�,.Љ�,��%��o���������sI�̔Bg�*̤��yڷ��U��� >�*Z\a\3k�?����V硿�oE�������M8���K�^��#�¥�]��v�`�:���m��Ya��휣�b�R^�i]wD���Y(-1��h"d�{m����5k�U�������Hw"'��7�`<��z������D�O������~>.����#�ﴞ�_�'�����!���F`۬�]1*�)(WIY-+B��2�rL/� ��c>�N�`��&��e\b!	�����ߥ�6�(�l\�v�tq��/���5���xe�*j��)�����p�^���Hs@L-ߐd��C�����
k�'m��]�[Y�^0VO�e@ *]~ ��5���"�	���)��j���Z-Pve$r��"c��Q��v����ޑg���)c~���p��|z�H��Y>|V�K>>nG�v�t�P��Q�T^�2�۶����
�1�/T C���f,��b�� Ib�Cq�Q�7��^�,�K��Z����if� 竳�FqX��S�*Z�,����c����҆<xSO�p>,grz���w?(܀H�
e�����[��|�["${����!r�Άƀv�be�W �-���������3gu$��/�j1`u��q��?����bE2�P� �f���Id��B):��N ����+�}�
k�6��f����v5>�靁H��@˫�9�P	���(�XB�Z!���[�jXJ<�]��`�Ѡ)�v���l,F��I�)��| ��@W�1j>c~���ys'��i��'�M6�9����?!0�C$�8E���D�(��a]X ;p���"�3�__m��`��3.]zO��£iJ#�^�C����΋��=�[���AyX��?+Zě��74��*���4�:�[G%�s�y���M��|��(�m�j�� aԞ=�4�0���r;�3��<��X�`TZ������L��m��@�{5Z^���Rؗ)�ԏ�l�ދgO�O�t��lE�y=��U2;y)�4���^5.^�%��,�G'&� �ٯ�Y8�s���/{�E(lp, �������F�뽇{
ʱ�s�㹅{�+�S�ˆ$��B(0����]�����|wr��,��~�v�=�'A���y�,���}����0�n�|�u��+�D�u���çQ*g!�Af?"}���)E8!$�W#����e;�T<ic���>�O+�N�uEX��F@��\�Z�E�4�ߌp���!��ЏӦ����9AO����(����8����/ �&������Kjg~�(�Mgo��R&�WҰ^��^m���S`�:�f�{|:ς@�-�{�.�D`�?�� �mF�������aB	z����Y1[��lG%�r�D��Z��0�@��:�[���[���M���:B��\n�7�l�N�i�}4���3�H��!��������߀�tm/�k|��Њv3䡜>/x���|U��A!f#��ku]��jas�F���������0Y�9�xZӁ���-�q_Ѫݑ��適>�ղ���l�#����O᎟d=��O=����i����y��B�>�ĪO��?�������<Uσ;�T	ݻ�+fg����mL4�@4��I���L� �3�d���
���2�#g���?a�Ⱦ_e�9���V�54��Q;yG��/j"�H�ajg+�՗�@�C�k�V�nuZ�f���_0����f7��4S�E��$�1q��e,��#�1�r�n�S]VV������I��`��O�Eu�:j�%�F.<�C}x�Զ���	s�r�5�oA����Q\�%��6Bh���wA-��l��� �8!�g$	�&��d�����X+�+����>S�xd@���\E~�Q������̡�#9R��}��������}�F?�NϞ	_�6�|EtȻG����[*fȸ�Z��J�l�+1�:-	��u��0�gB�hFT�@���kh��1{��Ay�7�(�'��Jz�������ձvLL�`�xTr�#}��|oMħ�zy�3Hu�O[�@SH=n��rq�E��m���Z^�2L�O��i8���zm��~M��Ѧk�D�/\��"���ˊ�A\��'��:��P�l
s�� '�^�n@�\9�>y�=p�+c�����r�cͼ���>b�Cp�mA�?���W��B"�J���>�5�p	����ȿR||��_��5�]�Fs��hÉ���A�!�RY�l����N���7	Mm2.������|��0K^��Ð`>�1.� �.�~�a�Zi�-��2���x{mJn�*�束�O��H_l� ���'A���E�v0���3W@�נ�׃!<t.�垺{b��ub.�W����ne��&�A��K	�9ϐi�$_U�C��c�� |2�\���Q�H�0�g�ΚC�J i5�DW���#�q�xᳲ�� ���zv=>Nh��c��ߕ�����j�4?�������-i-�I����d.�����Tc�dVa�w1~�=�9�:8��1=vM�l���(��x��1kroHA��p�#��mt��F�g���U�w	Ew�Yn�U�!����>j'h��r='롸N��mvlI�����k���:���Qu�å����d���{޶I����s��'�����S{����F?瞅���S�(=�bTV��.]A=I��n����YzV����|���2n�:�ѼQ�Y�&�#{UR*H�S�q������U<���-��@��-{ݬ"���v>y��fX(np��<���W�N�ko�CWK+-�E7F�H�ӂP�����+�[X1Ÿ��kd%�����SΨ��d�#WO~(��EΝ�?Z�oٌp�t�T#8�`3{�0�J�����d`Hq![=�<��r�!�+��W]�)eS-��;z�<��,TҼ,~���Ktg ��ڳ�o�+��J�Y]]��`�v?��*@��pU����ޟ�S�����4h$�Q�J%
E�ШdHi3��%)�$TN���쎐�:Bbۆb2O��Y�Y�:�߿���^�w��~����p߯�u��{����%��K�o��}ς���PͅKKP߇�b�XC�Jh,�J��a'M�S)��k7���J:�|�f&�O[��h����
�Do`E�%�Ⱥr"���y�u�ڮ�i�L���řV\K��H�E�dIC��4�1ִrW�Ps����9aM����{%�Y�]D��ޕMu�jY�[q�Խ ��]�;�m)�F��!�/�
��j#q#ٺ���Q��y�vXta��)���f]&#���É`�8�M__!�.ӌlxB�'o���\�ՖEtdІ5��N��ʝ�'���=�],v�tw���Hl�K*��t�ZD9���t�0�#(ԓ���ͦ�1��H�:� T��t���:���,OgJ�h�#�1��V%ئ�
�]+H!3/�������Gtb�:$t����ŘH�6���gf�4A��٦s�m`���R��:Y�]�ҧ_9gpVk���\-q�?�81����������#���w�%�C8�FS�PA�2Q�ѓ����R�k����&Ժ�LS�B����v��#؃͋�A$���1Ã�:��9_��^�g��k��<?_��I�Θ9x i�.�Y���+�9@g��Ϡ�x�(��3��$�&�v$>y@�I�!�e�fG�ڮV�%��IlN����W��O�C�Ğ'���?`h�Ǔ��z}+v�=�]��i��Zsf����[E�_�����b����3��
�Z�x�X�y��a�-Oi��jc�f�}m�tU�0�2���)��T�X�`1�v�s@Q�(:���XD|��@g/��y�j��"ZF0����/��C����G%��_�?dr~�$v�r1ֺ�a����&@�����`YR��ŏ��%��ʣ�=�6 2 zBm-NΆa#���H�e��,B]���W�g���I
'���.��'�b�Dg�k��e�/(*���ق�����8�Qq�V��ںM��)�,η����\v�����ӳS�.�������'d�X��+DP?ڸ<�jw^�,��S�>�A��c���i4�%�y�F��#��3a��	8�)lSU`m�3.(�,S1X�4���U[}���.�7y�>�̾�_���5��:��j���4dp ���Do5�[d�2F�c�"1�Vq�j�cdb�ٸ��
J�E¿�z���3�׍�3�z�1i0��]p�U2��q��H~S�B�B�w�G�"�
��*�{�?f��h#�������	���m8t
������M��0,xj^�<�e�#Rǯ��R*�qV��4B���]�[��l�:x�ʻ�Y�Q��y{�L�2�}��X�u�v�	���}'P�������@I=ϿɈL���O���Y
�(�<����M��C[�T�z�Lߊ���`��H�����DL�#�FFze�H�
�2���@Q�7���B�Io��!J�X��b��Iڴ��ӹ�Q/iS>Q�_�0��=Bh��i(�Pi��T+��#�i��~~~��*_����cۨ�w� �)9?�G��e(O���Rw�&:���=!���=qd<,�zx�2e�xł�2'O(�^�!׊��Ǔ楞��:� V������j���E��O�Ǒ��H��]�&�T���V������)���X�Q9J��-���ߝ���h'E��Wgo�J%� Ü�����y����%����8#�$��viT����y+!����rG��VA��I�E$��n��n�.�S;�&����Y*�x������ۙ��'���kb']��-t�J�
��~�%���7�˝�;��o4���Ź2՟�W��ؗ�L�����XG�|Mw�^w6oq(wP�K����(h�/_vOs������f����ʇOt<�y��l��t���ӵ�S�/+2ӧp��7+�/w1�z�/lMc�����}Ip���'� Ǫ�wH�5���>J|�蓶���5�Yo��㐡��t3�\��ʽRMK.�ǂ	e�m^�_}�7!�Us!Π�o�ܹ�f�f�P�:�f!����cT=P>��u([C:e����o:�2��;`U,�υ�+�^�ki�2��2���A���]�m�Apr;��>gǊ��+���ΰa؆��7������m�uO��������_HP��c��>�v��R`�o��l�C�����cLdz3Ф6r�8՝��-|.)����KX!ո0]����E�7N��-��=ޝ���P-�Kq�<����;+,�$b����ҁ�錓HE+ksH�������w��fd��$��˕'�?�ܫC�|S,���CNx�y���N�Ng)9��K�Kc���o�瀧���.�?�3լ��'��u����+����JNE�#A�x?##C����=�(�ؗ���w�~S��E�t�K}}=i.�?����c��1�� �GCV�e���_�������@��=E�(�m��/��h
�.�R�JZ6�	9̆�iCgg�OۂC+�B|}ۖ3����V�����X���1t�be�h���R���	%�ju��� ^t����`���ӵ^������9�.�Q����Yfn�&j�݇T��j�H{V���TL,�Q-M=�!s5�C-�����ɔ��<B�c�I�)�g'g$��1���o���k��	J]��<�l(9���C����6\���	�-l�z���>^��9�ӊM�/��%�=��lxD:����ṛ���կ,W�k�P�]�~���ٽ�=n�ߪ8��j���˛�w���\!U���Ef���2̚v�yυV1�[f�drQ����yv��u���̯��?w%�)��+�;����]���]���j�ΣL��Xyl���������i��xC0�\�]�]��&(��F>���x;0����qΏ��狘Umtx��`|�����Vg�@�B��y�)��ܼ�,�L���W�hP�Ӓ�?����s�Sا�� Ã���\�˝oFz�)(W�ǐ�-%�ۮ.'�}ؒ��_lE�$��=��|Y��*��oM�o/�`��+M��\'�'�w�W�@>�qt����ѽ�Qظ]N��a�=[�6���xԼ���>����P�X�0�5曆����v�w%1ӵ�{|�m�h+��o5!�_K��P)Ͱ�9��9�n� ���WY���pִ������YC���R���%ў����o6gM�L!����T�Pp[�����o������k�G#� l��:�j����n'�C����2���� �ڌ������8'f�L�Ȝ�f�r������{<F�r}�L��7�4���x�����9!��� #���BE(�ր�����辅��~ju@�%`�j�풙d|m���d�lS>���#s�m�fΥo���M93\�'ݍ���n�Si�֮/�%�&џ����Hִ����!oB�y���Q�zJxq5DvcP۴C��9ūq��7�t�>J�_����(����8H�ڸ�S�>y��H���������t�b��bF5Ѷf�R{�4v�_�K+��P|$Z�m�;ў>�f�]_8����X�f�1�IK�y2��}�>��*]�«��-�	W��:-`�M�Hv��F!��HS�&b�8%&Q�̪��[�pS�v�o6�l�\��ʜ�v����N�������C���BA��Y��#v��SY��⼇>�}pZqY�Q8�8��j��BKc)S�A��@��^�����]0�O��s��;���]�QNv�ei��)ĈY��ZϚan�꧓|�.՗�J�:wLĲ��	ɢ�?�q
z�"�[0��]��1g¢r�k�/0P ���4�fF��M���I:��WGQ�Yf�{ �mC�𯴡&A�CXE����GCv�.,&R4�<�1e�tљ��e�2������u>FN�	��WG/�a��򇶢����>^�>��y����`M�TmqP̊�n�W�q������?�1��;��v�	,L�~d�.sJ��(E ����5u�EQ�fY���i��:�`}\��T4C�c#���v��w����Œ�J�p�!(�q�c���Y!����Lm��e� "��$I$UXm�d���&$�@	�K�����c�<j��W�>��̌%�5�J��	 ���ӟ"e7��ƒ�;qХ4YԱ�㥯�P�@ˊ��)&�ksϱA�A�r�K��"�������@b��>F �O�����~3�)��9�`���ǗL�9��y�{�A2ω����~> ���k��m�
ʘ �m���BL��;�.šXsoddĂ@w �b����?�:=�ZeV|{�)���]K[.!��_���"܉}S	�B��`��*�G�X6�h%�����G(dv�y��N����9���u2�ξ)���=�6'�_P�	B39�׆��1����<�R����g���'�pS�
�;S^���[�+w���K'm}7��"&l�Ӽ��A�R�N� �v�X;u�l��֧(�#{�^,��5;�Q4��l�-$��x�sw��������]�>^�y����,��$�(O��9�ƿ��=F�K��Y%Sf�C3������$��e�{�W{8��im�}�p	���V/|�KK�ɓi��]qj�L�5���.#�5���|$%&s�=��C�1� ����Z~%�2O��+��$c�Z��i����s;�*�,�	B��rR[������KBii6۸4��8��)It[�(�4�F�;��&�5b�kh#M�3��(���wn�>lZW��?:D,X`�"�H#z:�|\���{S5�Ub����b;�����\]I5͝�װqF;e
�8Zg���X_�@��6;��HEWC�<2�(:������~�ߙ�KO�����yyy��"47�$���������0��[��[��Ry�h���F��
E��;�f�>����@�x�2���S�^�XJ '��`!�d�Sʚ�� ��ϋ6<��uo��)��J����u����6�K�o��-��%�����K>�$��}.�����o��-��%�߿d]Χ��d��8�k�,شtQ�k	�w��'?�9���NP����l��b��/�G���8�E�b��դO]���YS����I3�a������N��l��_��=w�=����_�����Ԅ��<�x�΢G�9�X�x���xYeŻ�p���lʷ��Lr�W���'��+�cC3Uߥu3� ��X��%⋞k�r0m���F����+�
�/o�Qx���H����=�0����Ig��I��Օ(D���u�'����3̓��ȋ�&o��}7uss�����L�n�1���ϒxmК�N�:l��������L�M��͇$Ѓm��.%��1~�;��Ï�S�u/�X9�<��kj'���5�r-�G�q�o�+**X��sx'N\O�u���fr�����|�����!�x���߾~}��X;���e����	�h�Փ��O<w�ɝ���>������!��XK���&�`����yy'���S�=_
�ք�������'��3�6�T�VR���/�?WH}nP���G�w�
�M�7|`ZC���hu����)\+#q��;�sVV[�f�]mt�'�����c��]�����KľL�q����޾w���n5��8�u���())��}l���>�����<��%�t&O���Ŗ��$��Dٽ+��s�c
��z۸F�]+�g	�0�����ݓ5�L�z2w��Sh�ME�*�՗s'����Z���m>��K�~���4U%��d�](E'�<����Ν����Y@��e�zI�K&����`�/x��X%��ܖxhZ�&/#����G���@�}_G�����/gg�E��1�8�v聘�ĜOn�x5U��[kIݲسg���7K���{�ʪ�P�j �h���ۄx��U�yRNJ��|֫�3rK˼���HI��K��+6OP
*��W���}IYY�>�٢;M�:�}�$��1�U��F@�͍����1#���l{�
�]���RZ �=�j�٪��u��a�����x����.��'$$�$���i3�6��"�����ay�w�=�<�#��t��|����P��P��5�p���YƑ/⍿��P�T��L"W��^�H�h��}�����¢d�]�=��t�Ѹr��"u-��K�
���N�
�	�]�FX����z�t:f�0�3yx�Ҽ��ɵ�����������W
��S2k\�򭶬�Mc�QV��t�o�uN�Hԇ�"��5	��ș qCR�����Ż�Yj�l�c֬Ys+�Ħ��� �`9�$�G^�g�2�Y�y}ʑ�	,� Iu8��j�+ٙ�����;�(��}��á�D���,z�֚彽�1�!����ew�0?|�p���=d��5�j�[Z���;1P�rQQ����_��"�R��h>�'�ؓ����g��QZVV������� Y�,�Nۯ��C�����E��x4�^�xx�9Ȅ�܉����x����v)H�7 O���d_y A�	5gq]��V�%T�-n�U v8�i��ݻw
�`�����H?	���e�4������ڊ�F�U�gj;;;���y������,�r�'D�ꙃ	N*�$I�l�䜳�@���TwVXX��E�~g �/�P�=f���C�s��ȓ�ʩ������ɰ��k��ҹ�o5����K��8�@���Y��\>����v�)l.�6ـ� ��l$"a�H�����>8!^�q�"�2���ֹ����꠨�"��و0���6�����[�D��kп�������UZ0e�jEp��Pҫ�4�*�77���;�(�����_o������&3D ���_�x�K��no�N����>H�J���)������V[FH:u�C����g�G^nt�����_�ǲ@Ą(��9�HBy���c�Zw�\i���颦I�y�!)���l�o�o)�eOw O��׸�e�p]�V�U'F�}����`u�h��j#h�8aE��\��I��
9A����~�@4�u��ȠT�AX<�a�?}}}e���5i(�ӭD
�Ҋ�XND��F��g�\q�;��?u�#Ȟ_ӧT�^��F�D�/O,vPШIZ�0$��XG:B��s���ψ���G�������\�Ȭ���Z�S8Jڎ�6
OĔ��p�3���3簦�8�����`_�l�$�����K=��K��Y����zezhl��� ^DP糳�S��?��z|>��
�����+㇓kX��<�Y@���T��c�����	3�F�ӹ�\�����dw?͇��SrEݜ�?)������X��X�|#��8 .H��.z���ϟ>�vR�%t�p�51�c�%�������s0���'���NЯ���Ќ	�Z����_�F[
O�6�a����0o����(i@n��H��Z�o	z9-6+s�/4S�U���l&(9���!�-_JN<���%H�6��
��Z��Ʒ�ՈWx08��Z�=�����	�����ju0����~��[|IFٖ��������|�>b����?%�>e	.�qV���>��V��Rɾ��Pv��̿�P�$� ��{&P<�d2&R��ƙ�!�(h�M7>"�=l��F�;�NG�1�"#�4+O������=_A��Z��KI��F��0z�\r)��V�t�^<ovtt|x�j��ϗ�9c/�:�Iݸ0�&-H\��SI<����j��ӳ�=]]\��IjD߲�]_�(��-�l�PeY�_����3�a-Mf��|(`��� ��<�{b��5
�q�[�)�9���<��]X$��HpǕ��ֺy�~!sI@A���_�&h_bz>D"C\C�za�����P�BfZF��cFF�6�#��8~i%?��}~����BHpH\k���˗焊'B "<�㡥�l2����u=z.��W����B0"W^k�����߲�ju=BGuʈ�|�߬A< �?P<�3���2]P�z+[�����U�m;���o�&:V�	e]�_[	�J���u�\,�E[ֳ2��4S�ѭ�����͑���D�e�SI^y�
Ƒ�e>h%��ڬ�0J�c�Z�٫x���0�[Éߕ�:q8�7��
�: ����ε3@?6-�hu��"�����X��y�p|����=�`��f�sX _�G���sQܐ�3ӎ\��O���5�m�v�@1�����7h��a'lE��`����Y4=h�C���	�$��P���Ȁ�%LTM"{��v�#��R��i�lBO���S���nd����c��pҘ�U��ЎL�M%g�h���� Z��v s~�\ �K�Q�O@ �m����J��@�/�<�qߴ�w�\n�Q�AS���|�o� �@����3}�RG@蜟�t �PCÉR%�A���N��p��Zm����D~P��x��6�0�X����$L����P߉��kyAb��SS����$$?w���E��-m�D ����ƴ8�Լ6�p/mQ9�b;��S� ­�ʪ�<��%��,eS�<���+��\4�301�<���f�!F�Ӏ��|��K;ہ��������G�Y�ś+a̡���'��$�SVvp8�l�� ��fNc?+##Î�7tP�1�pI�M����8��|X�q7��p�f8s��������1ϒ��o ��^^^Q � (ـ�,(���\%��m8z{��K�){{{;gg����b�yN�x��#vt,��U�|�! �K'�}�&�P'Z�PE1p�t*����u-GLjz����ȴz�'���T~��~���Qd ���|T��\N�-�̾Π%>�.k�d���5B�p%�A�b���<Fm�LiZ���\���5'�[�Ò�eAAA{F}x�S��C2�(-�$K�s����x��1	�7������gTy��
�4��F|��Y#��8`�����	�Y �g���sEX�j ����X��USR�K��Z�3��@q�z}P?ꛠ
e����e��_5�����j���L>�&�/P���[s�.�1捞6�w����ETDd"b��H�p[#
��䱱����p[,�@heq��+9g�8�UI�;Q��`pĆ�y���hsf����nNN���C�M��p�7>^�� �Ċ[Ʈ +;���L`Ts��MM�
�\�)��>yG�T�t�)�g�p��_��^K�t޸��y�>�tC�'x���֞#)%�IƝ����?Y9d����@��m��x�u8��V���Y��f6���ڞ�\"XsJ����%XM�f�!BΌ����?`l�Wu���(k5Z���'p�ף�f�&��!dw��[WX�BLG>�_r3���-?:D��!=�PE�e��w��������=���}۷����"�1�_~ �DSq&Y���:VHܴ�8��&t�F�y��g�-~d�%>��ضe��%��P�YXX����1=��?z
�)` ����BjY�tYY���hޣ�,�f�'�I,C� EFH�tΨ]FR�,/�b�D����͓��������3O�bWW/�
N}I�Kh�@q^b�&b)S������\mVP���Q��C���R��,/����]ڰ�����d��k��Czu��@PN2��8<KQ{�k:�O���0gB����|*\�/9��28��1n��MT�G�L�^� QU:�WUH�d@M>m���"͎���/��ֲ�xВ�ɏ8�GQd��gl�l�M���6O�t$7(B$)�?�VX<��_�I*q�'O�o.	+��&�Eo���q���#VA]Э{� 1=*��7���tz[��W-/y�% 吺H��#\�'Z=�<}]�f/R�)ݍᤴ]�.�1MnO%�8�+���9V�a}Z.6�k�__�H8��gh��Юh�#�:(�Qp�[�,��V�At[ �������}�
Tx%���豦��ka ���"V�5�^�SO0�J���9IV(��r���Ff;�<��K6:�&ЋU_�F���t>J
 wW��w�R��y3Pdځ�h5R�ǝqrrzO�l�4b�jM��.��[g�*"�"E�T�֊@��X�j9�N�q��2��Zq�j�	!wb
�c� m������<��K���p[&��j�� �yJ�r_���	����a�c\�P���#w�(#��8!iZ-��8���G���5>�Yپ_t��ĸ��xv�����Pe���Z��ə2�Q&�����[�?����{x�}�4�b��A+��C=h�C��`w(½���c�PW�����eQ���i��k�3�S�1���SS?Q�v�0!��oUD�2��yyy�'��o aXS��܃�e���4���Y�A�o�6���6���Ci'���;�##�j&�BB�c�;::��������^�)�-�ide�_ī�q�����6@��$K (�Q9߿U%eDEE����S'���M����42[���@���W.�����>2`ooo8�D��Z�/Xs�eJu~G�q]'䖖��s���x^~~~&��<����VWWǐ���(��	�[W�e���ͳ��/����8J=ej�/�A Pt%U����a��x�����J��$:��vǓ4�+��(a���S�œy�'z�	&9��� `�#ěڈg�!�Y���8	�!!!7�S@3��pg��	��ё`"@�&�~y��w��PHyrJ6���r��ǜ��B�ĨD�)){(<�6L��R����M-�Pϲ:�:,���b��U/�rw����ꉊ��Kӣ��'�j�~%"<(Z@:#�<L�.��#e�l�"n���h�9��[`,�Yl�ᘱ+C�w�v��c�qU�ZS/�a�I�s�.��?�k�iϞ��h��p�S��p�r�3��3��3><��F7Q���y�����.���!ƭ��_� �>�$w(C�B:�viA��Lv��rd)��������B��&����Ԡ�FQ���Tdd$���@�����X,���*a(�R$_���ܰ*y��4t��	����H>�r�Jf���mkKX^LLL���F��Jj��� ����	a�e8q�L�np�]g�?��`��.�o�}||0�1S�Sj=�t��8*! 	͉ll8�p]��L���|�O�ƃ�\��"������)D�IS�V��Q�>�ycw*΢���l+
��޽k���1#��J&Ҥd�1�'Nl��	B=����b�<�?�`u26>�Y�m�܅�x�:���<�	>�|�\龸p�_.��}vt��_�����/�Y�����}i���+^|8�W���T��{�$2<<gC��8�t�НOt�@�V8d�>�����[�Ŕ��^���?��p�9U
�[ww�a<���ד�Iii��N�H�w�*+QJQ��fy�'T&����f�l��f�A�6KrÆ���ʄh�Ș]L���29���"��f[AE��왭H�����$�u�)�2 6�>��{	6���%ǌ���-��(,$)�P3���144D�*�P��l�'�рqU���fnnNOy�2]K�!(����^�����e�C���'FRa%͖�2��Z��g��@{a`��šq��]���ߠ.Ȓ�T�݋'��ت�����o��}J�N�X�c`$�ܥ���
tk�H@������X�q��o$ZgS7���[F}P�Ћ�n�@�l����
�4�y:�]I	�ܓ���ʪ�	dޥ=�!�yU��u6��POS�hUU��E�%��~w�����v��b��u��l�0)��������Ap�^j[�/x^��<�Adt�X����y�v�eFHH�+����i�e�}� �Y�ٍ���;���*����("� � �
<���@!�.E8ST
g(����h����^YY��`0DvGiwrJ��|<*�s�ܘ���`��*咖���Rge�m���xg-�e=?�^*VR�p-c��ى�X��,���A	��0���̰���qn7J�S(�~Qeq�H ��@L�0����[�B��kEd��������* �����MފA���a8���;
�vy�`�VBBB�Zu�����zks�y
b��
��;)�q]�T���ɭ��t4�P���0�ɭK�:
[��$G���rѓ�[����B
=���(_���s�b��R���&3�(r_��h�A��o�⢿����Le
P&���5VVVw�\�}�H�c~/��u(�|VXX�	�&���@ſr�d��&M�UW#�@���"(	}���5���Ζ�~�/���dan���[�&��$�Y�%���=��f�T{��u}�� �Q�SX�S3NWRp����2Ț��3���G�[�D=i��z����75���T��F ��:��w���85㢂n��g�_h�ۏ��m�4��#��F�u�>J�&�x6d� �-���QY��Y����?��/?�`��|�-�"�iuP\�elMA@#��y�������&���/�ߓ��E�=��<��]���j&�ZB�GB���p^OO�~DO �/%%%ɓs�0;/���M e{SX�cF/b����ւ��B�Y*"**�Is�ޔй)����ၫ�s���6T�3~b�� n��_�G��N],Ėc�9��!іd�V@���>}�l�2u-��S�+���져�|�L!�����)�r�{zJe�x�;�7�<�Ig.�^Sb��␄8���F��q���h�ԭ������k�95� �S�11��Ȃ�@�k����LϿ��z�-]��MK���/�!$��������FAK�A-9eC���N��s�\��x�[j�s��A��{�6�� KB(N�SI̤�^p�'�?DS{{;V/�H*"�@�JC6u�?�6*I�9.��]Z��<kj�2j���͛'�a���F����,��o:f�p���\�
J���&M�uc}�<���R�-)i�8H��AW�A:�:�����Ɍt�*(ෞ����~|�J >:��6��ņ�ed���܉Ȋ�+yu��*C-�/C��?L�j͔��{	����r�^ ��k(7�4��$V=�	�U��ng��x�@qܤc�;���_�*�jkU��*jĐ������&L!�� )]��$+�E�?������p>�_]�p�����d���hˏ�]��㸮`��"u�����It��
���i��y8���f{�={���7$)���� 1Rx;B�6T[E�?Խ����STYY��8��i���kvv��^8��n��0X1��[�註�ɓ��H�ߒ6i.jř|6��5G�ʳ7/�OB��)�vv��ĩ���Y6�Kq������kɝ���p{944�:>>��q
�,Ζ4}�=cF��l���c��2Nx�������)������c%h���J�tj:Xt���^�s���� �3���>cFRYC��EM�hsNk~o=�M��RK�����"꨻:q�Zhd�_D�$vU�vu��
�-����dƜ�9��ܩ`c|g�P����:ܱ�����v݌2��@�(�;�R�[���}E;e���BB�ׯ�lE�!P���H2t���+�f�+��4*��胢�r�AH��������
s\��#,2kٲe-Ǖ����d�C��-	�v��t�רm���(	Md:T���čj����:w��T"��>n�JK-na�T��fM<�X��%,�V� ����iOi!�ˍ
�0����-B	d\�3��LF����1��G�\��eu`%����B�����.�P�M��8KV	]L�t�vnAa~����F��� �(��ʧn#䍠�,�~(R�=���fc��������"&�e��*��䯽T:�|l�+�*}98�h,z��Fc�*��E�;J~$N���[ϑ�-���f$u+,2�c�Us�m������P�Z~&y;�H������>��d	��ɘ��I�,C�QUPQ1DwlS�.S�����W[m��t�����I�f���Ѝ�j4fs�����86�v��딅E���F��`Km>|�ø�ĸ�A��u����d��Ý��;���b H���%]I�~`�)��,newi�Һ�e���~.Vl�NQG��� �R���n�����a'���DP���PE���� �&漁�???�-^T(>�#�uQ����;af�9�F����J��0&�:�!`~](�Ѹ;�Z,�e�>��m4�Z�`@:,3ĉ�j����P���� ���
��0Fe�??�I��j�o�����.��r��-,?����i���Q�n���|��.
rT���u�0�y����$h��ʔ�]��X����`��S�U��pm�S�P�� �hHS� �(�ni>���ゃa!���mSb���8�oKS���V��h�|��g�I-��dS�YJ-�������|F�����W����}q�f��uA`�S �A�������=�+9�2��`���F�F�����}H���H�ڈ���[Z>N���\��X!tQ3����ͱ��/씱
g\�-?�]RR�0�9�f�P���n� /��o�@9�~jRC-���0��F�E��F��<�e)Yp}��3NǺ�x�������f�jx��m��F���N��l֨����@{
JJn�p2�>�AB���#���b\�a���Z�b�Y���N�]�J��j�Lvs�]���W8��')��;-�s�]�~������ҌWb3��7t��y�A���r).��Z�mgt���$@�CЏ��{�pRL���!(555�������
�E��'�_��t���(�ۻwo����_H`��dd���h�q�f4���`��2gv��r`n?�Nof�s�љ�ϫ@G �W��N}�1ണ�cjr2�G\�ǣ��3���J����c�ݨ����JR�JY�7"ԸC?�ΏE)�9.�����\�����G�������e,5G���~*�M��CU� �
_gq^��E:)���w�Jbu�bG������ Nd�}�*��P.��>�4x�d"/��.�A1��F�V����W2~*#�E�E'G}H��<h�f�����d�k���erB��w�z�3e����e�{����}������p3�L���XRJ�WWYT�4w��|/�.����c�GL8t��h';� f//���˾rT���<qpwA�7r�����g��,��۱�����H�rRr��\=��0�1?�@L�����o�g5G����o�z��n͓��P ��W�but�Y9KT"K[<������S��#��������v�������>P,�� �78������s4�eTʍ�_m���,�_9G6t_΃���#��s �wU'z;2Rt��Hڛ��%$��֔3q�3���k��mB�}�l$B����K$���&��� �nnn�x��n�OhM���p�g��+W��%W�b�{r*G�#��S1{���[��w�U�┉���Q�эS�d���	0����?����P���H���G���P�&'�����Y46�?���,���.f��S1�@�����IM�y2T��b���@Y06�}R��ɓm1B��q9F���#�;�er�9�a����w˪݇CӘ
��C��1�l�N<;-�i��U��%���`����^^#sdM� �B Ta�s�����IU߂���<5o55I	�s���/��֠�F|�\��G��w�Śs(u���1%�I�'�F����	�(ऱ���`�J��P�Yvu�;|���	C+u͕5%߾Y��~i�@�!��# �L'�i��=������G��3Ô�jao�U>���S{���s.u��Mʺ�~�3Ф#��
���ohhPp�)-8�8���b���MT���ԥ����@������(��kMv��;枃��� ����a�Z��5�2�Y�zU��޼�Vi��P�37�[#e����9���L[�#�d�ɐ��S�ټ;���Y�c�����n2�"�� |�N����":RJ��p�Z�����_<{�i6k��ʷMv�R��8�8i b瞢Yk�x��
�b������Lf�=����,�_�?� d��k30�t����DmIKo��ĕ@#)����minc�㋠��N��P[H"�')Jk���L�	�bpP嫑p��1�oі�ѭ��wO��ߌ	C����������u�WJ؎���+u偑��Ē,vN�6\o��N5">����T������w6g�D~��Uw�טn�-���l��$Q�BX����.��(��luhv͊�oy
���Lg[a"�@�
�F�eg]�=�������1SH�Dtrtt�̃!�٪�*����-��E�����g6�N����\Y�#�g�:�!�RF����!�lLLLSY����m�;��"/o�u����������6������!PM�����H��<wvvVXF�kn�N�e��#����iH#���
Q���Q�ub2�:�
���3gC��a琒���ɭ��c���n���Q��bo`��m6��7�5Y�2,�N�
*H<��ġ[[��	O5l%6F+��}��U�N\�5�9K
����,��A�Ȯo
5D��x��0����k[�3�5@�q��\A�T���c�;P\}oP8 şξ�2#4%���(b�&�d�^'�P��i�L��
m?ť����-a%�iFH�?�� ��[�1�K��y����<�*,4t�G��N3��X]]]�@�Z�qR\������O�*_��n�ƞ���]��3��
]���ݨ�1�RI]��d��?}�*-)y�␻!0��3�N�U2�c#����Z�s	&9!׮]���	�C����s��ul�*���ɬ*�-��8����u˚��ZXvǾ:(�s����<1q��O��.gZZ�e���7�(~T~�qwԇ�sO�n���p<�>���(���q:�^c���ju�|n�FP�J��/���f<o*J�˶J����8:9�*|��BI�k�-1�p��0�Z�U��"Q#U�wGݠ�Z�ӈ~�m|x��*mL~�LG\��d���01.H��O�F�s[���~��VosW����i��|(���)�^�`��]�I�|x�]���szhx8����vŤ,�|w	mN�P����#p1�ݎ⪟v;�9νh�>|(���S�f�.q���zFF�>��F��H�&�r��O0S�� ���?}Z����۶m�ɰ����Ay�����f+�b��I��t�d)5:�� j���HQ��7� P0r�j��ǳ1Ϗb�׽*?�l��+d=ř2QlNA�:C����IV���qɞ?����)�?G_*�2]��<)�>�T��"�����U8[Ҽr��&�~S�a�w���u*pa�sNYD)���@�N�8�`啼�]��;g�-���^o�o��J rA|��K=P(0�U[���K�ۊ8�(S���'~�8%7\n�}��Y���R�0cU�ћ ǀq���ޭ�o�b=P[Gg�)��z���iiU	(W-���
i*�)��*����肂���U4�riiitC�xdVF�9ɽ��2+>7(�ڟu�c���]:uo6��x�ړ}c��o
6ų�[l�ɼ�|�w#�O7�/N\���xl8�|��ݛ��8������2�w���B�+V�)�M_�h���d/t_�(~������/_�|���;��x�L�;IjLl#���,}���;���MsR�tx:T��cN㥆�4��!>��}9d�c��)4?CΫtp_�n�JK�v��ƪ۶�k�%�U�.l��cF�3���vySs�/������nm�B�ۍ�eѝ�sr�V�}D������P�S�c�;G�ٜ���.o��~}�a$5fJnl:��ľ�z���W��]��۷:����Aj��j�W�����"y�ګg�B��i�9(�G���;����
a|{��!����o�������w�÷���u&����Zf9l��K��:7Z����[k��>�\ڄ1݅��ͷ��ހ�_�y'�}r�s����d��&2��@e�M��99���~5��ֽ}>6��oP��.5�	#��
���>�,�qv��<� ��3�U4��_fd��{[K�q]%�l`|��q��xX2��PoKR��,d�s&FF�I�S��m�@����aٹ��*����v��7�p�4'�=�|*b��cVR���Z���c�߾=	�9�A�@Z�,
�55߽{���uF	��ú_�\{������\{h����Ȉ���䋠ht�)�u�_3z=sTSr�����8���KS�g�svK����t��܀������!f��Qf ���y{_���ŋ��7\R���:�h8�|�ңŤ��<6�)<V�A�j�:e�r�	��~��e�aO�}$q�n��K��e]���#�ء�)�d�>D��D�G����IS �i��v'����a�z�PZ��QIA?�T��Ҡ%��w77�F�� 7�<������J�𲉿�a����`��d.��I&��K-�CG��d�M���N�={6fS����.�?���-If,��b������3��[-Q�$�Ӯ"l�KY�Cv�YY�J �_��j�"/��"��2�c��q	��wa���V��\��2	2L��6^���,&Iu��/������R�,N�O6b�ݦ�(���B�w���@��\l�J��f���Gƞ�.�����F1r���w�ܴx~�ڭޜc��taQQ'
��>��]㿀���@�-��O�Υ�����mD��V��o���S��c�B�̊�CSU�%%�$ �3rK��\�e����ߤ�Q3.�3jk>�60���%����}�;�ī�.DBo;�R�� �]RUq�rµ�ĩ��9��j����A�O]��'��J����0^�����2�2�+MvK@@8)�_�o�+!C�ގ�ᶸ�ޖR�HGo�-}�Tx��27���b/SRT'�rr�a�sw�Y⿛�8�4~Ǣ�oUI���ሓ����9��§�5�2�X �q�@���|FqW���(�yvuu�"{u��؛U��So��!��FJu� ��c�`��ħ�x���%/��0�܍��<x�`5�KC��杕[�Ғ�	{���������u��x�!_~�Ҏ+�4��U�sqI�k�P�$�3�CK ����}A�:��ó\?����գ*�+ �Nɬ�5�4coj{����|����8��CME����y0��A�JI���s�'�d��HI^^��#2wx�&;#A��zkC����2:R��]�I�|�ͨ��
��9}h�=aTϽ�7ⴃ��S�晑T��·1GpHt���1�m�>��[���G9��n�[e�<�� �q[�$�b%�d�޽���G���6�<H⤤8-:Y�m�Ɵ���&����q=�3J�SY�\���^���,�W
������I���
�	��\r�D���j�Ԍ��m�y��%$$�as��3:im�*�� <B2555姰=דz�������}�d�A|$0�c����~���e�ov�b��A�P8��4У~�(��2V-}���U��4�����'��*D�wp	�	 #Z�`�A��J����:�Pj����8ݠ���R�ۥ-d?�n�����nn#�E���a������p�ӄ?��}��m9UI�JJJeX(��X��ء&�ii[�Y��/8WX�ϝn9�W�\\}3��:{(zjrm�/S��ñedd��1�H���H�����TfM'Y�&f2}uu%C�[Fa$ �����N[��K�9�� '�(`6֟#�`�el���k�C$��5����dK��7��<�4@*�nR�v�^�����,�:����sa��j�-	�.��7ߎ���Ɣ�C�ݴ�K�X�!����	{��/�(�2�F�M�';7�S�&���26�7X�'��Jnnn��Ҵ̨�SD�	��訨���(�"i�Y���QE�k�=��ɺ��bbأ����(qY[[�'���d�j�vO&3�4��������b�!�8�b82DI�I�����S�֑���m�NF8�sv:+?m�u�L7z{�����0���D�$��pz�%Tj8!�)��ۓjg�υ���k�Ki))nz�D?����zl]<���M�	�XNS�R���d(�B�_��^wش��L�M�;$�����'r�{�p�ǀ���?cR�'�*��<�K%ۺ��[�(y�@���t��0��<גl����5'�����w�H�_cc#]?$-/{/[Q[[;L�)PwW 7�viW��Y��[i⵭��gT��:�A��/o�O�H�UA����	I?E������P���GZT´Q��V���(��W�Ț]F�'KSI�[�ƒ�����aJ��
�G��ނ~���9�����/�}����<���,�s�����̍���L��p��4�z����v��_�	Q��۫����_���� ;�{�s]J"��[+pwj�@\Q����x��ͷ��x��D���+o�ǿ���[.x��(�yak�1{O����(5־{`��1^���*�w`�ث��B*n��S+�w����$�OَʀΊ�I�-��������OlVB͉'w���ɚ���G/�2�����7G�#b�� ��g7�|N	(o�f#|B�x�dS5�lq�"��l���^"�ߒ}���G׭[���߭�b=y�u?� �4W(�O�nĳ�_ޯE�ree�E3�#k�M��d[��x�/�0��<`�4�^pkkkJZZ�	�BEQ��PR:�M�v�?z�A_W26𗯸�k�XK��O�>���=Y�q���(7�X���9�.�Q�NB�9E轛{"��Ӱ���\Ł>Cu;�㨑d�/��8�n)�0�U�W&Q(�F<�d�nR�$�
nfs��4����M���]]��� 4<��7��0PR+A�D�Q`�P.���Z2n�a�6^^^9����a�#����^�"����ߛs��3l����ب5ۼ�_�!���y�ga� � �~�b��4^��]%f��Ñv�n^�PD��.Ĝ���/J�����rq��c��Q�jR>I��A�+�mn	{z<�b��~d�b���X��]������ؽXzV������z�� d/�]��&�!����5�p�s�zn��U����'6�B�@�|�)h����p���+Zt���aX�nb�lsWD���-"��R���v�qb�V� ��v�?%;(���e�l��rA��Zy^ ���Cw��bܨ2	�f��f�"�~��Ͷ��)��+�I���{�����aL�Pn�O�6�s<(�Kł��kp�f�����v�oOyd[IP;��l�=۵1�M�¶u3��(	3.o=)t�#>��< �S�T�y��k���d�u&S�%�qHd/�n}������0�\�������瑧��*�e�B�.!�b��ح��?{^�5�T�����ͻb�y� }��É�Y؆��7���ěA�O�1��lq#B=��u�u����؅�3�=�Z���PUK4�]{�ڶm�7E�Q�r�XX��]x7`	e��G�5���5~+�e�
)l��^g�g"zI�Ph*�� ȟo�Z&(��p,�y���-h�孕3�psN����W4h������Ӎ.�Q�|�q#�3�>�X����"4=���<#(`D�������I��\��f<Oj�	E}�M��2	�5QUchV�-�VB�2G��ٚ5��~붉���~iI*�������`m�al�bD�-B���)w@f5Z�<�s)re�Xd�����V^�t/Gbב2�CO��7�F��6w���z^��
X8�*CU��CQ�z�A�]��>5!����铃W��F��"�~pJF�r$���ʾ�r�-Z��[v#�	��5=����
�=C��ODZᰤ��T�ķO�V��l��"�d+A_NBOV|��9�1c��{��En�=l�`j�g�A�/�rs���+�x	�^�GL��=x4Y ���/~RD[�эj�;�Q�ȝx&a�s?� ��D^�{%������� j���{L�<<bjU:��N��"{��M��������In`�cUUUx����^[[���H��ߔ�F�}$x%�{d؅˴���pD_��(�y�˯_�ЍS+� -���qy/
C�H�[��63�mnn��k�F��y�D�P_n;jR-�'��
� �ݸ;�yH�c�E#S�L�/<4��o1'��<y�2Q��C@
���M��0A��M6����F*"z|(��0X�p�r;b��8�yب�]�ty���M��
ٌz�G]H:��<>�H�&l�sIlZ�,��J��sm�q�,��7�ܪ�Y~�cj���`�{?�$���iy�,7�+~A!�0*%�e.6O��z��tLsGu��ː���Ti|���>�9}����rS�O.�l6)/����[�+ ��}�8m�]��xIA�K}��]�F�D�������(��h�'ZͫFPs|�"H>�Z�X���q�8Y>uC������C���(h�K�i�㘺��+���l?r;�>�P��$���+����;���]��������E%���]1|�}�T%�)ytd�l���/��C&t�&\.%�WM%�9׽@�ElS`���䖍>l�`��8l.$���ͩg���bc���Ԓ=Ӫ���G��`��-1(��T;:kh�M�� mT�i$�ȶ"�uu���&괪��l�x(co�d`��bȍ�Z�����|��`�?''��S�.c�4�\��1V��o�C��|�;s	e��IQY�x�����{� ��;���*��m�հ�sswI����f�C�[�9���+$�ʮ�V�ݺAA�0�q˘����,ǚt뢓߷"z}��ωcM{2z<*�ܭy����ȃ.��crjMTi���	O�v.�Gl�z��.���Z �w�WB�0�Kt���mgV�A�VF5ц���2	t<l�oA��Fnk:Wz��4[�o��F=D�͋�j.��a�=�ͥ��^W �s=��)z����!Yf�x>K:X>���D܎���P-}V��M�nz�J��eۅ����-AGQ'��Q��;g��o�v�Z ����ڸ�ǈk`�m�eQ��9�8e
w�)���^�F|�
��7s j__.�,�p�w'�����/i1D�I���̴���A(k�:��$�މ�D�Jx�sNl:���l���q�<tw��fQQ��Ρ�HT���=�sY���U�=f1���-���i�^��f���K�zNd�ǎ����62J����w���λ?$��Z[[�U��$#?����bS+H��?��3y� �d��d�qww���5�ޡ�-��2��@���#�5*Y�-~+�&ê(����phc�Ygo�>���B�Y�����5�(6١�
!@���x�Q���6��ˇ��ՉoI�u�w�ō��d�=�*v{$��B��h`� �1G���~Xo�_�˹�J��)���$�з^m6���`�]�ws�U��`�Q��\׍C���+sh��t��W���4Aa	����}�3@Y�~���zJ��4m���z<���)S��^ے}j>�Sa��YA>�s�ώ���R*��`���_�~����#��ΐcT0�"_籐����Hn�*���늖hH_Q��T��>z"�s��-S!!��QZ��4����������]B��Ԥ������3���=�-�������	b���á�
D�	�������@�Y� �5طg�Ac��f�U��x8�n�y��j%hFY�+ƞ�y8>0}kLOa3�P-��LP#S�3�8�;�*UR������)�rP���;� F�w�3���y2"�3��WG\�y3�����@y�P;ޕ��Xt�7&m�������N��"�a�}�C!��s��Bz�V��ړkQ?����1Q���OsA!�d3
_��*�&�ay+�V�@j�q�w9��E�.\�
X��/i�g�\ga~��c!�_�_�[�Ե%��������|�/E��)�[\u�1O�!k|�=�gI�����w�G�V6��555E�YQ�ZW:���qcwH���[_Ծt�v�"D���|�u6���?���N��!�"
����EW���A�}�{э	{���<R��th�� C�g`q0�6�I���&��h$~X(��7xi��}j����uttl���{f�ֲ�j�������$ԧ&��B	�I	�/�֓�>T;�a����ﴥ��jk�98?9Mi���	���{����5�}ſ<���8�m>���gyܲ(X��B�i	{Y/�!f��ϲ5G��wT�j�cE��=�n7Bf���[�94�����%,zt� �u�c����ϟ��v�X�����l�t0���誮��O�IAq��s����DeQҘ/}���h�(1�h��g���\�աR
@�:�DMd�o�@|���ؚ���3s
��\#��j`u�͏�6O~~���dSK�/w�\Ɉ^K����Yk���_�G���n�r��Pֽ��}f:#�<-�kW�(g�呁v�vH� �D���J�H��UE��u�5�M�����$ ��d4���$�c���$T�µ��k��7�t{�',��X>��Bs�A<�nY�������IJO'52C?+�C�i������v�/���t4���n%C��q�	֟K�c�褭<v��$�� ���(�݃���/.��)���zg^18ZQ��=�S#'����Z�4�s���k��$I��{Lq��8�C��z*�h_ߖ<��5�{<��]�*�؅/�sL3��,z��WJ��gc%OZ]א��&��"���\"��w�d1�PF��4�ou��	�������P �ʇx3��i�V�w-B�����.!�U#b��(������6QN�~�¹���Ѡ�V�� [�Ѿ�zw��k!�X�$��b��N�PaL��쉢��;�{Pz�r ��>��;lb�e�v	IC��~sL������OtjN���<�T�7:����浕�NCA~c�~Mь�?{�o�l�ӘAEC
�;��J�<��y�0����V��X;��_��}�2$8�`{��8q2����w���L��7��
Qhc%�]GB�is$��W>\��� ���R����ѫH��-:"<�`��%���+�m��r���C�M6��^�0ٚW��ϔI�F��Y�g%쏨�L���d��وi��5&��v_h����O�]��d|Muu:f�GҪ�א������Ʒo�y�N�"9���|�� �lR��ss`�����K=-Q���Y�:g�_woٽ�Tp�����+
�!����3b	m��:)��~fc`�`��'K���Bm{woQ��W\i�Ȋ���[��ͽ&ʥ:�����6��W�����4��;��e�ꛑ�}>%
A"/��uaL]�\Nm�*߼5����7o,���J�G�S"Y�����Ʌ1��2���z�C�E��\�iڸ�AUB�R�WP��=vS(�O�ݢ�5��� `����R��xr�����+�-g��<�&����c�h�[��Ѿ����g�
��X��p�:�+��v`D����
�S�ACeeecG�\<f�lQ��'�\���	R�{��+��oT��ن+�6�S�_W��w�/	?xv���􈶪�Y*<6�.O}�0��cA�f�R�_�M�J� ��9}�xw�������F���)��M��-@��4ukM�yd�H�w}o��p��[�����r�����w��6���,}=U��j�s;m���00������o1��
��M��aN�(�ns������Evo��^�*`����~++�����G"#�	c^$g�4|�P�^�W����V���!��n{_�c�]|8h8K&A"�T�	�1T&n����Qϊ��ʗI0%���k�RL��G��R������� �Z����nm�,w�a�3Ӌ��*�/���r�9���&�gL����&�tx�ܸ<��e�����<��2i(A�q�Q�D�衙�YײXm�sk>Vǩ�&W����q��Jl]E�o:���;~R�H�IE�Z�B`�6��J,�+���P}:όG�BcZ:�<r-̇(sY{P<DMvN�"E�R5�+��XE�����E����=ܻB?�t�U��0�p�`�h�h+w��.S�OG��ey9�뾚���<߁���~�
�!s,����(D�l"�=��Zg��=���
���G�3p��?@Ku����Rj���=_����^����L�8��k��^��i��/�Hw��(98я�G�t��
�|@�w��X@����s\�s�2/8R!QΨz��r��*	$ް�lM��ޚX����mn�c�Ѥ�O[��n��|ི���L=)p�����Z�-ᝣ7�~�:p��]��:��B����&�W}�;;]��R�Ie�xc�&�"��f*���lח�K"��[�U�C�t��{\��g�MGF�t��I��Z&�¥�|
[K�Ъ��x���K	9><���괟���P�d��y�����7*`
o��!ڷ�z̠P\�'�*�n�(�q���U*d��2���V�$��`c��3;�Wƞ���>f��z�p��n�b�E�j�O~��!��d��y�GW����}�St?-�j���u��_��̑���1�2I>����^ϓ>��*�J���]��d"���[��W�V?Z�Q>v~�Ґ��澚z��aa���>�
�:;��������Z[�k3����T;C'g��GcY�\E���1tsd�{	Ꝕe<�a��4+��e�|��-l�~�c�E����9(/�ۦYSZ��D��TE����X,�&�k,]�%>h��G��e���S�*1U5z���HcX�6P�u�v���T��]aU�q�4�,�-l���|�0��^־�7��~zW��{��ٍ.m��<�>�X>ͣ�j'k�*D���aG+�-u���&>��8�Gs���=�bt{k�4-��խ}����������B�x�c\
��9�iU�4��H�n���@]�=�N�h�5ED�����T��.�B��Nf[B�_^�kFPy��V�G������G�m������X'�Fcxa�}́�"�9�̺�Ci���(������s�Ѿ_���e,K�;�t�	�|% ��c�ij�*�cYn�n��*��\6��Y�k�UOKɤe58Ǘ����pVVV��W-"��#:21�{�v�dk�j���HgK"f�_��	��̶�����Vd��Zt���C�PA��1�|n���cc�49�\�kc!n� �i��K��b_�zf:��%D����iT���,�χ,���LB)��|J��<�pH�r\�	����8,�����x��H��Y�#!����A���g�L0ݩ;�.w�ws%b��6�����Bz<@O�H$	�c��yHp�]���hk��ЧbW�qow!��:�'r#�S�����p7�Myw4�1]ey1����j�鉪�K�i�FM#����i���=��8,i5�%�����kac�ϊ�h� ����ސ*1��_� �s�b���4M�Y��s���9�����ZK-o���P y�C��B	e{$�r����Q�'�E��l%n���8"��X�bUaв��[)�1��#亃��J8��d�P�J�S62w+������6V#��v\3r���ۅA�+R�.Yn/U���飏Wz�¸�o�%� ƹŬ�e^�]&���=��EV�
��i�j�c�$ �t�n�>�+X��ȿ� ׇ��,ӌ�	.Ó�G�0��J��!6t@�o@���A_��P�QOXE$kk�%ƒ��I�>���J.�MoszW�I!����:
d��m�v�r��$�a#6U�^L��y~q��xGEE���;��H�K{�1?{71�Cl���t�3p���T�.0_o��8&/�K?9������Ǉ��Ch�m�R�T���	���f_���lꝖ"���Ȏ�J��l�=�P$��-�����]�^��)��K5Q��8��w|x܄�R(�߸�@NJ�*���.I5��C�����o 5����k�Bs��H�=:2���	�:?���$���l���*F�D�&ʴ`���ÎR�c��<D� �-��[n��o��0��"p�_��1aaa֩�[�G�e��"S���u�
����+v?���}cIv]�V��["��U����ׁ%�d	
��A0m��Ph˾����i	�=m�����'�s�p�~@/b��)}U�� ����K��&K���*'i�q�.ʠ	 %n����������gʺ1B���{��U��L���^ z�ZeWd	�b{��`8�³W�l�Nt���?()C.��c����Jqs��+�}Q(��bbs8`jB��|g��P(��3n�r�A]T�)���$�I��".��"�|ZJ�s��]���E:�O�і�tT�Q�t�gx��.�Î�6��1�i���m�;����q�X�$��sQ�p�`���OGF��s�([�	�:7�ֈ�~] ��ĥ���v�����⟜�[C�Z4���X�/�T�J�+|0�޸[���Įԅ1!���Uօ�A)ѭB��EjXt֩�����-�W�g?�У�Ix��=EW�^u+����c?�%X��xB���IbQ����{�*�fi�fK#���GGG����X��WB�~WA��W�:��&ƜU��
@4����?Do�%���i������ɡ����.ז=�s�NT�
$?�L���n������w>��pOF��J1Ns��nb���9q�PfK�r*�aǋ*ҩV�#ցPt!UX\�SRbt��3���3�M$�L�n��
X10�����Ę���#� ڣ7��q�O��z#��߼R�[���<�T����5~�뚙6ڊ^�	����.h��z�VT�4�6<�e����g��nӿ���/\�rh�C���W��^r�����6��@e� ���B�D6c�z�0��(
Y�
���� pݬf/����Ry�a9�tr5c��>CJ���`o�6�ȐU?v�IL�Y��D�-A�&=WD� M��Q�pU)r�{�{

!��#�;���[7dN���mX��S�A�H��r���}Aľh!����
�;K�4���~2��	9��N7Q�vD>t����g�ea>�!�Έ��E'~"�x�>h��,u�h(1*ڂ3#�x^�r6�u�0�'�U��{�4�)"�Qߝ�tk��H��W_����� ֓�5�U��g��K�+�_4c���_�Ah�(1�V'��]UG��}����&!�gS��N<���@/��І���R���b��S��aJ��"�h�M�[`�6�s�*�{V$Je����tH�Җ	dC2dT��cnj�2���8�H��os���x�$�9GN��Kl��𢡊B���C��R �x��0׃�4F��u�)���mH�~��e��m��|�y��	�*��>YFF+�6>H��-��N�/����~+$ǵ��x��f��Py�ڏi�5ȄBTr�t�.�p@1� l�NY����\�9�'�h��m�22^�u�y�U�^��*D<.�6�\�Q���c�i�<��&x�Ω��gMT��\�p�V# ��;L_AQ��؎�4�C�5j�K}���U����=;�A��H��+���T����v���>�gBm+J����^�d�ᎇ�������.·���`�}��#��m�M(��92�"\,;K逎�!��̙�'�k�I�׻5Fn��bTݲ��D��"�iz���z�L�-�9�rfF����~�
�S�<b����=��Z��<�4�T����[�-���DT�3B(����K��.m����|�\
j����0�\`��t�������C�Aa��>�+�6/��,4^�����*��� ���}��}d;&�����xJ�ء.-�sx�.B��N(�~#U�>���}�a}���x�7g"Bh���+S&��P�Χa�{�\�w#۬A����Xc[����X445'O���>:��j�4h�A�D]J�E�	=%ƅ��t�{D��]m`W<_��K|��-�<�I�u*��.1�C��)x�Ia���Ȝ��Bn^�6`�je�x�N��r;���\����"�	�1��_�⓵�kZ4?!".S��
L��h3D�⓬TcbD)��N�YY�"Q<�D��AwM��A2j���J7eKbX$"ǋ��Ί�>�D��V�v���(=���d�P���o�նP^��ߘ��zd\�⏅���n���^�6����緺if�Y��,�/5M$̭|S�.�V�<�H^ؐKd��c�hր��c��((s� \��S�EWƌGi��7H����FP���]�Z��Hc,J!c���WD�y�nm�X���o*E��6LH� ����]u�qˑN�5=�i��'����Z��w	φ|��
oK8�v�$�[��7�_��C��2�;Q[u�
i�	8<����b���ⲝ���Q��v�n9�6�K(��\>���(���Ǭ������;h�ӡT��00�[<�t.�C�P�s�l�ǀ�(��.;��.�.ׂ�f��P��F�_K,a�W���Z����gx;����3�O-!Rl�ݑ��@X�k��L7���Sj��:^"W<�.��A_oŬM���u�S_���I�E{�vI�IyI�����3�I�C��.�-H��R'��/��誧>猎�J�f�ڌ��X�|�)ڛjb&�"�zJǼ�Tm��8"�$6{��E�g$�a___7h1(� Em~�6Qlh�-\v��ǌ��� �ֹ�!n@0��D����B��Rï�0�Z� 34�+J4q�.��s���GjJ���7��6�`}�Ay�>���	;�����^�ʶ��%��bE��&��p�|����J����r�|�܁�*^)We6�!� W��i�S���������/ ��9���I��:���:E� cu=�}�2�;E7��2��/8��PTB_���r)@[����y/����H�vA�6�u��8GnБ�$�5,=m��� ��P�M|��܋�a>��ȗ�d��`!�
���i+�C����z���!���>������R���Ĉ�e	��e,���Q��@\\\Q
�N, .LI���r5ǒ�?h�N����/?�6�5�������glb��p� pp`��;� ��~Ӓ)��/k՜�I���\4J1+��t�>���->C�6�x��qq�3qy�ձ,�GP�Ğ�/?}F䳔O����赎Od��>P>��p�d�E�-i"��t��W��D��7q3sWL��4�
J����S���H0�Y�����RL�FzĻz��P�9�-Xh��sҷ2�L�a}��r$��(����o@�t$:}vVe��v3��̚$����6wn�Z#�Us�����S��bz9�b��rԉ]H�`^C�������n�I\� ez��
����Es���E��3�Ǐ����I��nb�1(��'�W�:4�Q���2��5��5(W5����}���K�	�gn�"ӡ���gj�f
�rW;���ئXˎ+)����@]{�>I�=a=oh��sà��~���D���k�Q��et�&��'M�����ܷHj��߼Ÿ�7�z
�qLIŜV�8��d��f�F����!/�'�v�x�0�9V:�n�0�(y���(R��N_z��i�:7qziV�Eņ;E�D���F�SP���)g���(y�O��ys���;Ґ�= 3��V�a�����26is�J�11ty�٪�NvNl�S��w�	eV����J4x[[������Q�kj[D���}B��T�^v���Z����f�_i{%:�dj�(���,T��D*c�n�{�Vs ��߀s�q& �ɻS:�*��B��iuy_�!3r���Շ��_�^rqZV$+Ж\����7un��M ��@�����E��G��VhE[��-�q\VQ�=[EE���I���������4�d�i�|
ǯ E�sp"M*LzXn6��l߄l�_4��Li��.0�'��_,;�<��7z�ƚ�{�"�f}rFg��F'�/~��" }w��>-%�Y�慽u�9�A����6<�� k~o$/c�:t�@Y��zеԏ5ۉ˪���R]�ۍ�����[�l<I\t{٨V��{3.n��"8���"�d�Q���������$�4��)����%�)��i��z���Y���ϯb�4���+��I���k�JWĺ/p
�X��m��>���3s�XdY��s�"���xן������/��ײ�b律ⴵ&� ��ZB[��_7[��ˉ�'���Q??��������d/(�u�,{{���R�(BHӽaB^GN.�T�������-X�P����Ai���0��6�D�ӭG�dH~�Lfʇ%J��䛬D����`��`�KVQ�w��;��|y�������L�u��1�9��P��P������䀹i[���-s��S����I��������y���C��e.K�tkϓ#"��.�՜O�x���I����]��KPbӜ���#GrCo��.��@�H�~\cZ�� *)Ɩ,��-����^���:sI؟q�UQ��d
�V/�����c�M�V�tc������jv�}��r_�c��Vp��ag�-C�&%?낌�2ΞQחQ4|BD?F�s��ζY.���K?�x��~�$	�MZ�I˧?�I�Fm��y�����Ͷ-�z����\l/�ԁj�J���7�jS�7��_C�F��4�d��֒!��ۜ]?�������|J�5w��A��Ľ���nH 4��/3������ ���	h?/�X?��q�y[�g1�s���+�b���\��R]� �p�_3S4�����|�`��6Y�/�Vp�K��~d+�]O����'�|�VW�d����=×�DU����>G
Y��d�tYsb�I	�OO�V�I4B1�QJ�"߂����}�)����� ��b!����1�/v��"4�3T����dn�7`��"T��kj��ͧ�6dY�V�N�鿇(h�Z���a��P�#���N{��&�X��lL̝�izw��^���g�т5I]���r)P���j�EJ�{8q���O��{���i�Ґ��Ldg�L�!��z9���3I�S�͡�!�Lm���+�V��C��/�zsǩ��H�n���xr��W�44�Ox!���c���P�4�7w�N0�	բ����l#�?��+�[�]������r�:HVXۮ'q��j��#�:���F�����Q�ݽ��g.���8�~)i�Mԅ���{.Od�	�F��ͮ/�� $�
��Z����Cd����I��v�՘�d�P.Rq�n`�����9y���-b!���L�Q2�𬍫7��z�&XL�lҢ���͛-j-s��TfNaaaZ��?]���\�;��VZ����=\��b@d��[���[��O{6p&�3|DJ�$��'C���o��c�8��E\�*-j�}ٶ^�7�)Z�k:�]��G�"{�bּR�6]�w�%�e�F@�~��ږ#�k={e^{��M佃�]�O��b��ݍ���G���xKP����]e�n?�D�v�J-�G*��H޿���C�'��	��F�&kE�wT���5�Q��ӱ�]�Hjz6�<6�ҁHT[/0;�5'����')�i3�ޛDQ��0���i ���"�p��\R�ս1��=a,#�eVw���+�ߑE�U7)�6�Ns.�1M���y��&g�ScHݟxm^�v"�囧c����1�W_�;q���I7�秤 �e�0�. ��!��̀,Ϩo/()�<��o�@$u5��e�=�L��[������3��"������5��hTD���T���[�#���b��R.�6�}����܇C�d*���y2�S�f�b}��F^��g&�_Ify�\���Ə��b�a/(��͏�m�3X�qN��h��w�9?�z+r��$�T�l�&y��ȘP�`ˎ�#�7�Uo�����^��Z= �3�%�ۥ��ѣ�T�H�;��~�M0���?gL���#I5mK�
�h}�c��+�ε�w/������kg��'��h@����h�VE��jW�B���X*9���6̹�^�E^]�GMH5�k���r�<Sg�BRS����\>V5� =������͊���͙
�%�S��������y��EÚ�����4<îs^�sB�;�O]b�i��#����tΌ$կn�����Z��8�39C��\1QrV�F�&���(�D5�	F�̇�{<�I@luK{��RpD���d�C(m��1@��jD5�zq!��q�
wD�~,]U�+���w~Ո�R{�9jο3�3F^�G��_��S	�׌<�T��_*�9W1ƍK�t�l#.���3�%S���]���äΥϳtJ��+�ڟ�fA�9��.��ƶ=�X��a[��b�0��.��1icZv�=4'U��,�&MΪ�\5�����T$iX��齦�II^~�:��	��?�4����������n�܎�JY狐���E������ ��'�_m�)ɓ_�@�&��!��A�w����Zh�m�TzB)\J'EL�*-k"'��ɽ�������kH���(���j���<�'mZ0\oh���?��lI4�����s��&p�O�K�鄅|aW_~�:$�B��=Yfz��c�W{�z&(�݃\妡���c��v�֘��HA�M�E���݊JI��ʧp��f �C��j�z��GoN0��$y���2e_���w�r_(�:�`M���^~��q��u|u�����.���2�;d�v8���D: ��\| pV�x�=qm���'[[�LC��E�Y�ԓ�����9WI�������|�������1��Qf�}�s�1�M��W�B~��n����y��>O�W��{c�h��f"���"=�$U�J��76=`�ѱ�^^<���7���K�jo��p��N���@j_%��R/a����ݤ:�w��=y�ş��;�-��h�F�0��� ^^=i�W� <��_OZlE����Ɠz�o�ym����ɚ�X�o�o�U�u:�E��*�j����2���[v������h&Y�br;}�K��a�?�.�F��F�<)��ꆚOUj�
�T��F`�G��b�X�'RIqX���䥟w���z������|�ΗG��� Vhc8-vo)Y��R�P�C� �Ԏ�����������Tְ�Z�ɢ��e=!,S|��g��|5%��t��c�fr��(������9�?�*���dpKs�4��_R��F>��z|2�2Պ��ɾV���G�����!��m�:����0�C�򷏯���[��,-�W{��垭IQ��ꬨRM�D�wW��6�i����mq_�o[����\30`rt���.��"G��$��w6xl��&�������?a.�,Rk0���Z���)�r|�ț�H�"���5��C��̀��/?���l�GY�al�u?t�=4s��W���7����?B\��'%�D䔶�,$�Ψ��ۘ%��0�"�f�C�P<��~VG��F7������*��oE@��>M��q��R��mR���E\~�Q\ET���q�����`C���RSW���>S ͹#����<59z��#^�e���ڒ���2�SXJK"�6�9L��|=����hH��3�k��%���\^m�>Q��RF�&ҕդ���~?	!���k�?�H�(���/��x¿�mˋ;������ |o�U**���?>���A����nw�s\a���������f ��u�Tqc�����	0�U��Py��6F���Z���ړ�"��R�%�Q����׃���))� >��:��_����A2����n��u��E��|6�����f�.y�����E�ʿ�-�$=V\cmRJA:�U>x:�bɘ�\��UZ�T
ō��;� ޤ%ݸ�<���i*BR�bJ��-�'q���l]d*��;�5C[�D����$�C�ҁ+�o���&�0�1�M򿙙�b�!��8ȝ�_Sd5���^X���)���8���^K�k6����Yb�;7tU3o���Q��1�G����b�i�@��.Ss�`��*���f�B(����>�mX�8M��-r�����,�c6�}���*��MXwJ����9x��7�� � ��7j"�Ú���st��P*n9�B&6�)s8� ��ǧ��
�\]T�%�16f����S�7=����lT�L��h���m�y��ƩfΔ#��U�%�lip�)�S'���o��9��y�����)�z���0-ȥ�W)��[�ѷ2���9ØB!{��t*�HϺ$M��zu�Cv6��=֨����{��J�`c��f�,�'�u|o��6dFv;�y>�5 8�O�-���6=���؋������=�6Rn[#�R��ߥ��t���Ly���7v����=3�9�g��,]�@u4�d�t
��4�g?��K��
Ƚ����?|�P{�
DnD�� U*���0������!ޑX�֪�-�"�v�o�Sy{��B�p�fE��_��K*)����� hej�l���}t���:��j�]����C7��w ���@ͥ��Y fRf��3Mv�K�;[�M	c��6&O��4zaa-�%-��Ĕ^�B�?��N��<cH3�,���'ͼ �������u�b��pE\�����ƺ�����,���|�v�IGn"-xV+h�&�s�.�&Ś,t�B�������L��v@m���o���'��U�oN����~�*�����$}��@�:��7"#�v�����q4q��0.L!�ܖ���tNZ���YI|�̣�PԒ6�����w�}��ݚy�yC1�w/� mP�ܓ�;)��ܙ���t�ӫ���� <+�@�bm<��^sZ8{l('�,��sڧ�p����1a���Q)�踁�-*��K-��,��R��2��b�,h¬��`rAH	��[�ҙ���3�-8���	@߫
!�Q�uv�T����j����B�-�$l5�]GN�$����A���&=s���VD���)wܥ�8���q�;��X
��E����ωEĥ���@Mo!��m9I��1Y��$t�b�o�����E�M�al;P��C";���� U�C�:��|��pa�HB���0��FM=�l ����jF�u�uZ�,��vi���p�9��0�����%z�����4�3��`O��P��g��zL����Qt&�ET�Ĭ2TN*d�I��Y?��	�b!��ͭCW(�K�0��Z-�����~� ֲdyV�:����V(�|�%�~��V8��If�y����������S,�����`�����?M��~0��d$���a� ��4-�9y&���=4a�}N �(d������Nv�^����b�C���񎬟����������	�\���vkŜ������H�Ǆ�=�����~�9�Sh;�V��J����&j?_a��8�Ø�% E��(��`YP��B}L^�NEg&�nc�V��Q\m�R�ŷT���	���E�?����L�(�>L{���R��΄������+m�6���d��ɦ�<dz����Fؐk��
�^��������s�:�Ҟ�+0���z��d-��n�n�Ie��*e�
�K���u$m����.� �q���^7&�����#Y��I\��Z!L��u�5cL�/��]̝��<� ��wi�H}e
e��n��_��+�%!)��[� ��dٍ�SF��Gɿ�9o.�>��c$|٭!/S��]�F��*vC�JI�	�صk�VQS��*����HܸS�p�|oBߨN�P�M.����p�fj����Z����3DP��0����ʓ�w�U��#��V�����B�%�G��+*���,
οπ�O���G%�A^j�׋vb6�H�/9���k}��jna�њ)�9��./#c�5��&M\Lt���96g�QaJ
L��%�^��!8�龘ZB�g���GB�%�9�{��κ�Hբ���8ti��%A�|9=�<��>s�6�ן� 6M�ⴲD���s`�YQ�����c�^��dOk��v�i���&_�OnZ�.SrbᦹFލ�$']��Al�@!���ǡ���봜������FV�'��������0/�w��"o����ڼyϳW|M��5s8m[��ɾPen諔�(&�K;i4L4��L�,������J~���M6��i�֧����}�Y�3�dV1 o���u����]!q�� �j.Tg=���=��d��p���g���1w���?NhU�l�����ќ�L�H����ڌ4�kϡˁ&��7�B�s8�@O��ّFޯ��:� =�-���:�z�$ɼ\��d��D_���B�Ml��%�r�'{�ԣfL�
�Y���K��NHRc#�2�ˡ���0����xtm朖����H�l~�|���p���IQ�r"S���N"�A~���i���oa�8�qz���p�͌���]fZ��1��.���d��gn���)d��Xa\ߤe��&a�L��"A�փFB �[�sda{�k����uЈ q`eG��VM���FQ�Fu��C�b��Έ�VFZή�bw_����e��M�"��e�;PZ�E��j�}��+�'W�-�J��
b1�[5#oK=�,#��*������+1�jzV�G����}��O��,+�%3���fŞu�����1ov���x�x�8p�������nV>��Q7#��89����]cX?eSw}��F�/��l�er']N�\�m������r�	B�7�F��q:EW��͛�]o���06�*Rb��,��iz��=_ZG�G�ٕ���N�޹�Ĝ�I�^�5�(l�a, rK�ø.����о�FZt��j��;%��p���]�ts�27nt�,����
V����:�m��*����F�@,]7����}u�����j;�]���m׆��Ɉrl�QU�����O����o]T
6�j�49Wd6;�Q�J�?�.{�Ű�+�Sjˠ �/�/��?&j,&��W����6i�E���s�X�ŀ�9sg<����S�Ӂ�����F���/���Qc��v��R���}�����g#�8tk�$����f��8"�r@�>'<��;�u�@pC�@�^�
�K�ls�(����$������M�,T��ϰ�zϲ�ȇ��L���ƀ;b���%�g��Y���f�]��[Q�-��1�U�EQL6��(�թfU���T���\kdb��ͻ���LS(J)5�w���J���n����6M!�=��w�#Y����j����^��?�:J�a7���e0�m�H����{�R�����f��;S*���ef�����?��	���75 s�x_c�ݯ���>�G�;Oy#��|F��j�lf�{�ύ���puˉd\�lSwǋ��I�����"RF�/6�F��ps|��d��#i��H��-���DGq�����Q�JN%�L;�S����ڔ�%ǣ�+,6��:���w	��E������?R`����%�c�uĀ��+N6�4��9�T�������7�V�_5Vo>,"���2�ߘ�N�������"�SQ\��N�MV�LrG��/�Ͳ"WS䂀+���by/�T��=;��Ks��m����t�-6z���7?�e$�����/���>E_�k������5���}j@�������A߉E=�X'����j2442�I��I##����a#�<-<M���l��F���'g&�F Q������O.Pi�^�)Mut�A��޾L(_�kV���ylyF�qi���<=-�O�R�/�U)&F�����$u��x��Ɣ,����0��R�v#��CϘ���`�xJщ.��RO_��N��V 0���2��dY��Vj�ڥ��������+��j���R�ȭPYn�'d*S�.�[�R�&���=���P��ص�cOc��dP_Y����e,��93����?^�s���|>�����<�9g2_W�2CB�l8�o �]��b|�9�zŠZ;�'�hͻj/���3�~��^[ ��N��.B���Y6b��̥|�8�S���&ùd
U\�%��bE�D*�c���M?֏ B�X��)-�0���M�Ȭ��;�ڙT�J�d"7����jޯ��S]�w1�GG:���)?�2]�*��������`I@�лf���+[�<��B)���ܢ����Q�r^+j"�𷠹Xm���(��$!�+bI)������(j�k���46w�_�B��A��r�\d�q��Q?&�s �6��n��D4��Q�Ws)1��X'򤨅�+�
8t�[ӫ�SXb���������@UX'5�w0C�p�G А�ZE*F�������a]� ������^��q��p�.���	����6o��D[B�m�掉Y���k���5�z0uM���9eG��H�a��l���ޥ��j����a���'do�R?_���˾T ��韜{�OV���TM%C�(���x�ݰ6�$Ѓ�Z{��8�(�>�ܨ�Li��jP��[}�r�Pڸ���;/�,]��>Fn��
��?����_"��
H�f��?_�~*Ew�fFa�1����L�U�8���I�R=R�1@k������S�׹�?J
Lj-G�������������Z�:���FB�0� ������2TZ�փ�i���s��.KͿ.%fS��\~ig�\� �[���n�Yx��$�3��m�& ��D&C\M����f��|�)wZ;�a�Y\:/����ї��f�x�X�+�i����B����N�z��1{ �_���w�8��0�ެ�#�A�L��g����.�տ4j�oٔ1�u>��|���ɧ�e�?�kdeK	i��֪Ň���0%礴V��P��Ai�:rQ�?��hX-YC~�
Z4b�����2�)	o+(i��|��a�e0�<]��c}U�8o��\c>Wؼ ��oh�t �|�	���O)Fc3瀫�}+���,C�V���]�6pV�Tc�E2o���a�֭Y�$�t���/�l����'�ᗀ�S��ѶoX5Av�����ǒ᪷���?�\�� �F�j5���3r�!����"�#V<�\c�����X�\�gN]�V� ���s�����tpV��Ӫ�%�\շ��[N���(t쿙A,A�y�h>,֣��*4��1
�?����!$-3����xP�~a~�&΢��#����pb��q��3�N��f�����9}��<��DKA��(��]\j�����!��ak�]BL^�z ����CQ9SCg^���<�7�J�H�=��|4��,��d��� ��7�գ�Μ�y�u�J?1�`L�M��=&_F�2����\TV���Z�\Yˀ��A��j�9��9e�"8[�Y �D�M���f��`�:}Z��Wr|lq�$)���s2�φ@�n,���R�$N,sѓ�@�4e�E�??����*
|r*G_mīڇ���꒙�t��	���M���<�ɪ�f�jf��&��Cq�z,#M�0cMd0��P�%�4i���O�	�A+á���@����O�0�@����gA�}�������Z��s�a�$k�'��vJ~c���rݵ����DK�|�]v����d�� ��@���9[�"�0��S�|=�. ˑZ�pM��(szq�.�F:�\�&2��EZR�-�,���$�?H�SǀS�"�M�\��6��!�)�E��5a�L0���u��t�įP6F�
=bw�� �m0�~�-���ڧZ8���v0��w������@i��~z��se���J=Ȇ������, T_җd���Ϝ�MцCndH��#�Cm�V��)�>��dU`x&��{G���g/��E3�f3�D�$�9xڬ���F�Zm貦.O���	�b}
3�km@`��DG[�$x���#$����y�P�E�[8��Z�_�|��b���-
��`}1ZC���aH<������F3�Y�_W^<��rȚ�JK���m?��6�_%_��6��Q,w`o��l���6b�x�:�y(�G�2�q�U�l��u$����|�:Փ�Ű �(��U��$NS��+���]��N�XNX�k��9�d�a�=}���tvB%6C߰�B��0`�9lr��#-��[�b����x�(#g����=�m����k����s�/!��9 p��t'��d�7-�2�6j�!���
�#{5��ĕe����O�G?��4Aƥ޶pF�߲r�3�9�E_���@A��0c�-����(��=����oQ�ɩwJ�{+y'yAAJ�Z�Yz�~��K@�@���{fЄ=&g���3�~��Ф�\5��uk���h�G©>Y'�Ճ�=?&��)�D���.�(-�{�Y�? �2�`����k�3�q��Dӟ��|vs�gx�)|l�� } ��������-]7��,G��G܇�MY ;r�l��כhEb|;�b�\����)!��jKoZ��O?�u(9`�o���w�J{��_���La���CO�r�g���뫺9m�� ���K ���|d�ˈȴ���}����4�ǋ�vEU�FNj�U}S$9�(����Yf��v�_$Y�&����2c�׭?�/ k���:�{�K�k��S	�H��=	�8�w���B  �h����b���'M�*YK}U�B)����z̆�	4@�#Q�M \}�r�غ�]�W��!-�ӥ?9i�	\Gn���s%�X�M�}RV���6#	�)��0�X��Db�M�eΠ�*��� ��xr�����ksx�id�����K�j��;���Aw�i�=��9����^�7+��ٖț��Ҷ#����P�3��B��?_~��4X�;��k�H��D@�q �� �:�UVN �a�M�23�6IS35����ֆ���W��%���\���
�V�Y� �Z��YN���Y�!�l��쫵��D���[@�-V!��H)�J��YZ۷V-��ؐ3l��̩���V�,4�P������0�C>�Ӿ	��$`#wP=�cy���
�-��۰���澯wҦ�?9�S$����p���%jb�У�K�Z�͋����G�{�r�g#X�d!�7��$0�D���KK��]����7�,�� ��<��O]�>�p�`��.9q~e�L�+)��B��O��z�����>${�ݪ��rĦ�}�:�iZ��X5"fK��2�n�oWz^h�Ð�t�
v+��	��9C�{��Z	��	6�/����7:϶d�BGc1'�p.݄Ο�n�]�[���*?A�dx�����8�LT�@<��i����f��H_������$rIx�1��k��Vh��#�<�@��{�8��}�����(S�qp?�(ѕÒJb��}sף�F�8&��E`B>
�i�^1�K���a����S�?8���t�u2�M��"�z@�_�� j7,n�t����$�t)Rq��9";�2��[;Y#����i``��^�<g�R�2K��	�<�y
K�G�E��u��~� ��i��61u��:�v���ם�r�D��[��/l� ����b���+�'���d�n���}H��1)FTׁ��<�FQ?{��i�����g0����� y��f���pW��<�P_C,(_7�·�SY����\���	�{q�}X�
����!�kabͺ���v s�Ь. \�ՙn+�kJ����
���;1��X�vԎ��\�M�4�`?�El�wW-(:��T�?A"�m�������6�ΐ��.�{�y^��d�$m)<���bV�n�����W�t������#R�
zu����,��,���1ޕu0��l[@d4=�h����z���P�i��e)���;G��at��^[m��cW�kq��mZ^蝄�<b��t����\4�G�y�Z��b������*uy[�Y��?K�DS"���P�eM��>.��oV�Ꙁ+�H��i*��@��ϔ=��B�q��<��I�v֗��:g-��y*���U[k>�.�V��̑�]��U{X�> ϱw�.~��ŗ�2����E�.N��Jv\���(��5mn�T?	��b`�&D P����Ta�Ȕ��^��Z8DՂ����^��ΡT����:3LxG��g���Y�~SB�P
��p1��w�sL���i��5�> ����J��/QM}������Mln�-������o��b��D���������Җۄ���J1�91�&/�S
�Y�·[;���j+����C���t�cz� S���.�����Q�%|�z�@WV��~C�œ��!NC��0�GY!�C^��_K�a�]�� ��*��J�3�R)>=�,>�s��a��6��f��ne��0G��(�^� Xc3��Hb=��Nd?��+��"�Z��Sr2���ć�q,xB�!���38�.�R-I�-(���g��4_*R���S�����Ю[��=K$p���eBa�)7�\(n���o�i���hi^�ILN�)@>��z��~k�2�����U/B�4�@.�'��˖8��$]���� �PIt���V�9���~������NΊ�LU��I[*�SN�K��N�C �j��N h#f�FL�Edi9���ޥ
˨:�@��ҭ�j�fj�S���B.����6��ץul������b��76x��r��P~.zL���A+ٛ���/e�_�U�綱p����\9V�Ҝ���4�m'\�%u����'���!o/j\����ÿoy���^My��G_d8h;�o���-���"ʚ8����'�&T�&�MI��9��`�ޡ�%ʸт�S��>��bE��;�C>����1�d2V�=.|4�-f�\� &�xʕ$��D�N|�����*�zj��?l`�~�Z��EȜi�/�� '^�;H��Eќ��/�UZ���7S�S�����{�ظh���Q�����˫1��}���K\��?�,�:*eM��!-R�%�nW2[�!���������B��T�yl� -��e�-��m��瑚Ѷ�UCh�
�3&�Cv~W�E_���ު񱓸��cp��.É�� �b��r�}�,�V�7�~WYխNei�]��ӣ:�lI&�X�J������ǵmЇ��;A��<�.��Q����Yd�:�
�%3��m@�yCغ7��㧱��2��lCC���R`V�w����BB�9�􀇗χ�`���՞�g=��kxn}᪤|t�Y����dAvI���g�ݮ�*h��
�7�>X$�3ະ8P��vi��(�LK�����ھ���W\F8��p�Np#��AwC��sĴ��j����q�I�E��:z�>����FHb�n�GS��y�E�R�t�J����O���Zb����p�Y ��o�7՟���yr�p 8�)�p�$��3���N�a�~z?����K�-��������x�w��V������񌚼�.����f����PK�X* ��0jwA��b��
M�C�J������3ป�*.�Y0oY@�u�٠�4��$X���G'��Y{(⋢:p��3%�^��Nf�v�z�P��A��"�l'lE�;��Jē��|s)��\��9n���_f^$zs�G,߽d�hR�9$�3��Ch���-���-�����gb�a�K�eee���d��ץd`��[�I;��`� �}O� ��HFx{f��\�\-'���k�佷�x��0^�#�ֆB�vtt\���v�x�4�W���F\���j���k"HST�	���\M$���~��vq�+%w?[a��d��%V9w(m;B��/�Q9D���YfU$yi�eX���hP$è����ג⊊�fX$��V:Û򂮜����<P�
�,G�/`q	|�̟��~X�,�JL��rA��چ������J|b
m��H�e���t ��K���?��6��~�K���3�@+)��f��%��G�C{�A���$sd�]f�%]JJ�R�SOi��q�ȇq�!��qP�i�_���ȼ��h���88���-28��z�6b���+�XB �ўJ��͒>�w1��e����q� 7�wZ�e��)P+STTb�����Ҕ� ��.쬝΢0�߈qUڝ�2r ���Ӏ�]��@	�l��\��~�,��k�M�;7db�kZZZػҟ�.Nld+�3r �Y�_�R��>� ��ޗҳ>i���V��Va�1D�E0�kϭ��a�����EC� 4���DE�A#奂v�J�a�ڤ�U�3����x�К"���rに�srk͈����y�P�aH}k3π��S��
���{E'��t��_C�Q�g]9�\J`��G�ť��lL����r%,�9U�����͏����U�M�]��#�1܆ϓ�8���6�:�FM���@�Ȧ��K���>��7,��?Ö�,�1��[OU+VN�)?�$p.�q,��U������P�����,�9�������:��E)�N[��=�K�|��C��uL#,�����z�f� ]�PФI�0�']�ʹ�e�g��z=;�ٸ��Z QhB/i���<{����������hd��0����9�����*辪�j�ӏ�|1���Ɗ��T��� �k�Mi�z9]K��}πG�RR7�	�㭹����ˮC3��άUY�%� ��)���;ef]b�?���2	�����6A�����>*%+�֍�j|�y��Hܣ>)�3�Pf%��JSo�~T� <�=W���j,`�Q��� "E��(˅8�`bb��3޶w��J�6���c`��^?^�);qV`]�;���M�p"�� ��[��@���ʡ!{~�;	�:�/l�{䇟�[�Z���Es=_���{�=�րᯏ�zP?�SA��d�*�>��"[�7�^��%=�<D���k�������"� �[��%�Ƭb[�,�7��U~s
�P2K9[}V�wƛ���+�6�M���+2�|��M�ڵoƊ��4K����IY��X�P�|���Cc|m\��2��5Rzn<1�/:_�(A�AN����K5�r���z�#e��b���\Ȉ�]�fK����a)ω�iLi�Iݦ�Ȩ����Y����n��4?��U�5d���N�W��UĞ��&'�p�+��D�GC� ��q
i�%F���ٰ�z6�'���B5�Ĺ5��W�3԰�,h�w��e�c~'�����"_1��.�'�����	�
�^к��c��d����OQ)Y��sb"��7�Ŏ7���Sn� $���e�yVh���IÔL�����(8l,w��X�ΗF��u
���q@NG�w!�g����l�z��^O�3�{c�<�N}�e!�U"�nZ� �giK��1Il:o��3K���Ok�=C�آ~¼ҾT�8f�:�M�(z�mL�� ��bJ$�$u�`��M���Q�g�k���2�g[��6�ǥ�2��p��[���%&����w~�B{=�&-��N��f���Y�m��s��$a������x]����(z	_���jϙ�:����BM��-n�I��#�G�`�6�z ��f��؜������(��.��1 ���Ng䅣�3G�D��A���'1��Ǔ�'���
iU�YJO@Z�נ�*��,�X.�MR����=6�f/o]P���8K,;�����H���=87ϓ�48��d3�
�\Z��V�E��<���Ѡ.����5SWF�՛�ڋ���oa6ܨ������ނ�ٮ�M���?E��Oʭ��0{o��:A(�O�*[���7_��,X��DȧB�w`H�K�R7ΰ�����m�f�ΐFjir_h��w��.�����=���TjZ���%�)�)١�����kJ]|=v$�"�t�.�B���(�d6�q�ɦ�0�'_��[�X�����k	��S1��n}W�X�֐���>��ڑ�W6��K!H�x�N��|��̰�jf����q�C�`����w8vSQ1]��+J4����:�^� @B��xX�>�O��8,B
89�nS;i���k8V~���[P�GGG�0��Č��a�E�<b=h�$���>E1$�%[��s�S�v���}q�5��܈�J�R�ܐ���$��e"H�-Ѵ�5�!�~����*}~��F��(9RӔ%���!��.�VT)`��_�V�����/I�7�b��a@�;o�?V���<���������l�Ѥm�1&�~`idd$�*iP&�E�cAJ�����U�<����� �`��tZ���z�U�8�Ջ^����/�=�	<˩x��T3 ��N�k���G�^�_kB{z�h�FD ����~��,���A[̈́s��J죀YX�pa�Z���U���d�N-l½a݆���7$�B��'v$����x�!��Hn�If>���Xgs��%o}��"p� �,2=5��s���s�%�)�#�rW��Q�����z��)�b�Y��>x>Z)��7G�y{F�ft��złA���BP2bޒY���& ����@���$Y��r�	���V|��F�n%��B��t��$@#��#-���0���v�?=��c*q7S��=��qR���O ��n�X��ϮZ
 8/���j�k�`��!���Ub�:�ښ��TOϜ��+���SF�.���.�a��(H���+�~�9M�7�Y�BMRRU3�Dce�>�RRcaշ/��봣����N�r4,���D���><�l#��9�Ÿ�]�4���T˘����
y{��T��>���/Q]���F�-B.B�NSKl�DP��`C� �ч@l��ǳGǹ��}��齾3zL����{��>E�}q�,53��y"���3\=���������x�A�}c��?�k{�s�ob�f����
'�#�%���b��7㑟�^>!��PS�j4|^d���Ic�J�@�x�L�����<�0���j�Q��5��^`H�MQ&��4�!����O���"�ow��4���q�e��m=�aV���W��$z��<�.&�UJ"iOVti�/�����8?�1�2�4�j�jW[��lDr�䀈`�1�/���&9%3IX�
簫�X��i�Y�qx��G����.�y`��g�{S�e�
Jr�5�>�#�җ�NƜ��2���'�
�(�u�;d�~����m�ˌ�b�	]}�!� ��t�ϗ9�9�gv28���Jf�r�����c�O���}u蠗t��!3^KH�os0?��*���Z���H�&=9tUFx��mUxj����j��j����kϮ¬����>�)@����Ƅ�s&+XL]�K��Ģ�\ϒ�F�ӏB
@�bN��Y�#e�pR��I'(��fr	ܛ�K��[yثT����d��}�lِ�O�x����3��;����888(�q���^�5��(*Z{�.Q��L��v�������F��@N؁f���\�%�|*v.���rD}�PɌfPH�{�Z�+��,��і�>���Ȱ�mmmOa�3�ᦑ����IGE,8�B�a��c&�ډՂ�:�\�H.�{F��%l�K\O�+���d��ؓ�Q�T�q���SlI����A�!ۤ�u,�"�˓Wr�;�a�^�,H��M�U(��ݰ��:�����F7>���&��ʿ@��L9
j;vBK����͢�cW�|��	���{�_�y��̜=pc��� �8���8o����%�`�f��{�����a܌�T�P�&�u?{����cb];�	�J,�X�����$��	��iry��.+*)�Sҽ�֠Rŉ���DX�7��pQ�J��$(a�-�r�>Q9�o�K��o�����BAk͵�� ���9��~Mj��R�D�S�4����ˬ����G��R��6)� ���5�����ƛ3����`<�V�u<3i,�ڵ�"خ�.�
��-��>W�ڤ�6ň&G�M	�g�M?�C~�U/I����Gy"웽۔i�;��wן�L���Tg+��A������UMu������f/�dH䣝��~�lE�9����d������I��ڧ�N�*�|�;[=c!J��x���	E'*PG��U�}���C%������k�%���j�)#e�SUS�x���y��Cu��'� . �0��;�fĥt���Z|����oR�mU��C��7"H��
X�exݞئ�J7��H����}G�᳣��a>�h��WD���i�@�����@�ދ�	x����kg2c�n���6�q���
z�������n���5?�wǙ�ҍX���W��V)��z�՘
,
���%�U��:���`fcס�l9a�j�5T`?
�W��+R�%�K �N��(]Wr�*W�]�Ӳ�<7�E�Ԝ������ �)�		eNa?�h����M6G��k}� ��n��pn�u��x:-o��ްc���B�d�Uw/�`�'�>#H��Wb�sJT穽sssE111j]���l���ۤղP�'}��������4`�,��{߬7���+m�<u�1��T��q���VH�?jP�̯�;z@�%E~f �V�+-��G���^�zT8��Drf�O��sF���'�D�Ϡ�߻<�}Ɨ&t5��x�I:Y�/�^綆>2�8�;4�i��ſ{����P͝l�\�(�˅�/%�� �
pA<�����p���&j�x��˫�!��&J�q���.o��.t,]Xdu�?�w�*h��Q�[�����3[�N���a��w�w�sm���ܴH�k���4fc����9��Їq��1�S׀㚺��|� s��\BdK<_I̟��F?��r8u?8@.��]]�3����
ٌf��<���ޘ
�k����,�߼�ؙ�}[�e�G��ӗ���B�h��!ޛ���eH���;~R�9�%#A��|[�&q,j�~yр���w�|J�� ��������2
��bJ�u��;���>��=?�{	�oW����
������^�o���G����08K4}M|���UPo �J�נ!cA��g׺Oչ�h��-��|���B�Qܓ�ځ���i������vx��m��I���*f|��D?1W~�W@5�vdr(jW1�E�=�k��s71�` ���D��D�|E��P��d����Q�$�j)�+ӗ�?ÚN>�:�,��H�<��v�w��.N,�H������Z��V�
yNOѽ�z��S�Ntc��x0@<H�J&%wYsEtf2��ۅ����dK�
)!^W�����	^�PF;�?�׳U=���m؏g��v�5�w�|A�����1d�*R_U����<�c8;�vCl�ގ�\�����o�H,M�`ŭH ��RF����:�N�!8reen����;sd/.���a�J�v%��� �w`,>�e�����y�Z�����@�G����N�H�2��Gy�(�
�!��Eu���e���3��0�.@SR���@������Fg��N*���$���}HO%|��W�NʜQc�� )����Ǐ�V�HZ�#�QO�1I��A�� M�M�O*�Y6��?VH��G�Jb� Z_�(J��'����n��G
[� 3/�j����;+	!�
[��B֟�:�%�}U��
�l3�f�*�(�|x�̋�Ê�y^A���'��P�?!�xy�(߁#}ԅ�2-D��c�X����$�>��r!��~ N�҇O�C@x�C�xͿ�g<ƀ�2K�x>�骽�(Yܹ�>��gb�^Y���0Ot6eWm�gس��u��잛\J��@M�1���
�M��д��*.�Uz�@�;Н��ff��pZw26�g�7���[��1�SR���j|B&������/��p"��*������//�g���x�K�+*sK�b{�y8NI)F����W�7��c�v��� н*�u�����r/`tw��;(2���hVkԩ|m��>�?��>E-��<�> �F�Qi�|�
v@�w���P6%2�B����;Mps���N�h���%Ǭ��r�ĆX<�#����\:�𽦀����='�ۄ��~0>E�Ja.�D�W���7��J8������G޲=@�wZjs���N_E�!bC^p��<�5J�L&S�{ei{@H�	�"�*��٫,�KX����h��Ő��̰_�M�Gu��>��1�)��NQ<PNޠ�c�"��y�xuwbt�UP3�ٔ\ӟ	�u C���0�ί[��i�����Rk���Z{�4������G��J��w�~:�f�����%.N$a����l���B$_�,�	XF��	Y�R`����(�� Wq���_�ʡ�K7!��N!����Sv�O�H�]�%,����`�&�xx�����F�B�(Ȅ4)���~��f�A˿Ïa��5ԷCP�S��2P�2`�Yj� ����G��j"�jR�|�ry)�\�"àEA*�,��
�} �����*S �*o�bO��� ��c����\[�߇!ͰS>�,�J�����W��Id�i��u^GH
^��?���$�m����4�՘�斸��N��k���!�5�m��'��81���Q?>4$��p�`��:��6�*!l}7�Qz��t����R����8��9�Y�P[�o�[Y9&I끯g�F�ID�_�SO w7͘������%�p\��!n�=>)���M�L��%�� >����C�����������Ѡ�������(��_��R@��3��r#;FC�gi�#
��P���o�}�j��"R%ol=�Qi��H!<&0ï������I..�h�CH )�֛��c�r��CJ=�luM.	��D�C�l�OL���,����Qw `P�.�ߧ�\v�5?��j?`����E�@�~���O~�ɲ�v4߽��֜eӆI�c��9,�A�7�G�������ܐ���S�Г8���OcE���ܹ��>� #������FA�� �QT���!g�D/h��Z�%�|6�9��6ZYA����K�����X5^���s�>���E׆�C�ۻ�A5�{�m�M:�W^R<:����8�����hE%dz&�%=��B���v2u3�i�TGa�9t"�;��4�L
��4V^�mA=d��п>�cA9t���N���2)��&�|L���y�.T��il[�����t�G1|�����5,]���s��x��b�!�sӻY�Dg��O�!d��E���!��o�烾vJ؆~��f���6ĝ:w�'�n���!����N��@^iL�&���UYޮ�E�/�*΢�ubo��n��Q���H�fd�t2!�8��������4L�.�V�xR����YEI�B.��8��C~3`�̾����R���RD��0�E�sֳ����y�Ri��Xj�mwOO����J�gC�@�؇��}�������i��_������f�׾~£�a����(����q3	� �z�1�l��J;x՞"{�o?1Qv�w�����	�+��8rs�n��+���5Un���M7!k���!<^���ċ��V�t1���,��YB9t�%>�D<|"OPG��s4Z(�PNC�PZ�;1��k��bib�߾�%�f2�����UI����Z[ZZ�:\� �:��4qK�V�-9RZ ��&,�;wN�|�����{�*�bBi�ӳ�=vt.��Sn�Jn_��F���M3N�1��
쏅=�T�����g�������v��u��Z�J�9%�p���	$�c���\������;|o����F���jY[[��?�^���fjb�pʫ*�{E���o��옷g����Y�'���O�.����}��0� �8�t����ɬ�X17��&��Q�,���R((�ɑ����O��eeKx$?4	�W���E;��{��pM��xm?�\����:��>�we܌�*�x��VVO��T0�	8y���\qbbbe.�o�> >��
��I'�;|�[�$�X0ϩ��k��z\JX(�ap�D���M�[��V��jqtҭ�oC��]K����������j��R��D%�4�À�sp`�א�7��\d�]SWw��j�%+�ؕ�q/Y0O	A�HP������OԷǥ���I�Hz�%��5�h���*~L�=�!�,�A��}�;~U���W�?m�
�����)�@��x_ �?=�-!E����'!6JY^A2�	���dX�R��!$��nD�O����a���}��0����ƃf�@Sj��x0Qk}5�QB��%j3kN1�R^\}�"�I�p`�� �*�@\��'���_��-)ᩘKo��$4` ; @&p���.�z��(��@���{���-�7�j���+:���ÇUٽpڜ�M�֜��`�N�-�j���d�Pj8� ��`�/��a̯�&�������fC"���J(w����������*y-����d�'�}y����@}��������7��ڡB���X��'*jI!80h���9�3�l���*��?@���K��*�q>~��0]�ꓭO�w	��΄7J�7<?���eO;����@��)Vu��m߫�[@����NS��U��;�4���%��.9%nO��)��&O2>����j�_�� ��]>�ܕ�M��T�q1����
�$�V �&�Ŝݞ����_<�;�;�)����jN+���M��7z���.N��V~P��哛Vs� %g�#J\���IpI�2�;�֎t��Z��-v;��}	>s��l�nHopXs�_�#�/�~)�����,or�'����m8鋟Y�i�����������y�ж��{�5��?�Nw�Q����-���h�v�p�_�Q��@�M��c��?��Pt+��\��������c�
�/i)ߍ���٥;�&������SJ/�MR�t	�7�WV����s��:��+pf���K��.�8_������|lg0�m����к�_-�7|�R�&�:�ۖ^+�TmSK=���H~��������\\�n+�Y���ĕ}LL;��S�t���]����L1���&V�hM`y�oʙQ�Wb�>˿�Nr��PcS�) ���]�)��s>�&.D���	�����i�.�Ja�4xݸ�Z�۷��o�O������ŷ��ʦܮG�>��0*�U�^g��a��n�:t�6(xk؁b�*�p��z��%��`�2��B���u-}��ZnzyW���O�5o����~��H*���N�s[��C��	
�ޝ�^�뵁���|��p��R������y��Z��o��w4&:z��䭖4�f�<hʣ�'�ݼW��[Fz�餯I����'�!=uHW��[I�c�g�mBI-����b&�/o�4����r�w%�q���w3����t�[`�⎬n��%�VH��N��J�{Y���O��6VD�(@z\���b�f��ү��o��K����@�F�����y8aSgI������R|��)�`�s��G���8�yr��y�9'��t�6���N�Mu^ʅ��;;�k�TYBm����vu���/V�oQ�D"�V��<�P2��4q����io���/-����þ�9���v��w��yn�̬�T�s4K�s���|]g��j��Э�;'�w�0�<Vz��)H7h���/��35��j�de�ZU�/�v8�o�w{$4b%/��i�;ׂyYd��+G:��y��碯��|#}�%�G`���w�v���<V2N���2����Mccc�U.�HV�W�k߱���{��T}�gaч��Q�kd쳯��K�-�����}�RK1�"����XA�D��q������N����|�tb��ܴW������9
�yTn�X���J�q��
k��@�?�pN����;l�h0�M�V��uv'�hQY�>�?�X��iz��%��?m}Bm���}"iT�����\��Y���2��Ƌ�'X������{1�Ҭ��fh��*�y��%�^XYYI}��G4���AX�랿�k;�Z�5޴ggx텈���r:�g�%�1-�e�r+��ǥ����h]xF*�]�4<�.+''�^�������ź�+�������L�W�K����+ߜ������>K�^+���h]���Ja �rr����<-sAeȁ�r���*m��XX�8���}n��%�F9`��c]�l����9�>�3���d2��VV��m� ����׾�nv���o^�M$�0��ٽ�r�L��Y����� �(�Fɱ9��	�륍�����5�=H%E��$ge�|�k��?�; doǏ�1����{�,��ݹs����>n���l5��󵶳��Sͪ����/�)?��>`y)�2~6�{��/�|V"_$��A�r׎)��P��am�yQ�7ͺjTq�䗄�A�w%���@��f��S��!=�N���B-�om�6n~&��Qf��k�w���;�Vs�� ��k����n���@���ҡ|R��o��{����_��]]������E�M�qi}���cx�]}�q[��� ���t��o��쾛���M �\��v�����`dd��������[䵛{}d�o�w���k��Φ�@��]�\c;�>�(TZu�]�j�O{���B�fE���M��7�#^��>�X�qǍNM9�z��������g�o��J�o,H�< w�색�j�b�B�%��P|Kw�gC���B�����	�RI�a�#�<_n���<���"��I�F���\\!�����5]�!�f�|nTh[���-96�Na��nUUT4�v��I�l���p���L%�l�����o�H�i�R�p;��oGt����F��v��wX �[z��'�_z�����)�G`��P?��i�X�x�j��v�f��U̥ٽ����uY�rRT@����V��\,]�t�]�qO�Y\Z(����n49��x�>/�7��y��0E�z�ݟ�?�-��0�~��]x����)@�q�Ϯ���vT8�]W����,�$�84���㲒�^y�h�6kI�ke�p�;o���#���a�4���k�Q�ht�����eSDˆ.����x��G��&�u��B7�P{��,&�[�B���0xpCCdܠ��B��w���#�ϥ�Hy4ix����Z�<옱��?�ˤj@A��GU�@��mHgxvtekG,�^Z�J����DO���׽��`�^F/�$^�T���A�۷�b�M��P5�ɰ���.������
�'�2~�Q<g�b���j�j��]��mz��|�KL7��0��Iކ�
oo<>7�X rɻ=I���{>��W��M���a����T�x��5����j��c0��ݝh $7z������_�-h~l���$];JU��q���6��"d�߁�;ݸ��}t���ڏ02�����O}Q��/���kl'%�;2�1��.F�w!���)��4�`���{aӞ����~�xg�.����`A��ۧ����:lJU��"����B-Л�k�p8�䉮=��ɋD��+r�x.���o���S�\��=���>G�Z��?���@�T�MP��;��]�m�?h�73H�~|����Ŷ�J���Ax�R����N;���7� ��_����r���c��zdjjb�<���a�X�Z�v���I)��{k��e�A#��3!&�
b�l���(���;R@@�`~����9�R �M���J�wנ�
�2�:���:?�N��%�S_�u��9|����U}�����>JL$v��4}��A��c��j�~}c��Yug�ȁ
0�~͵Ϧ�3��_�
cFGh��d�=<<*F�&����휦|�Q��e�[E��ϴ�Z.�*xʼw�����<�s�״�}V:^�D��s�I��'����`�"h-fp��{��c\��O4P���eL���D]�M�*��NM;����]>p����HOʣ~1��nĉ��W���]�J� �@��~�T��7�&P�?��E��͕)ߘ�y�V���A�c�r��#���U'�\CAѮ�^c������Ai��{����@����*@��_� �m��nRD�î�6IZWIX�yE��s�b�Z[U����@O��T�C`R.� � #�|�F�BDg��c���EGs��� ����������~P�&{{{#1�9�@�x�|wbk�m>iӞa��"ݠ)�r%���I�a���-X���4��;�Oϛ��͸�-�8a��3D����|���Lk��X��R։����\MMM?&��$eBr��$][���3bo����d�_-//�z�f�-��ǻ�{���e��K)���|�"\�H���\���5<��� )7n1>�ip��Ӷ�e�1
0��,�䭥����=���ǺUz����D4�v⻤ݜ�Z�	�B=��ȱ�1ء��i)=���(�0��UC�U��C�3���k�����56�"��*s:��+����m�`���EwF�����Ǘg�+W0t�h���E�=��C)����7�N�5>ǧREs��,;4~I��O�TI1y���tM�~����e���G�����%�T�m��P�H2�
�� T2mlIi24)2�d�2l��D���XGE		�mI�2��L�6Ŧ��?k��������w��:�w=�}�ϻ޵��^-BZR�A�LTD�mS;zyМ&,_�)L )�bHQD��I�;�Z�L�
��I�o�ԓ#��}��d�3�([8Jg|Qa~)���3��S��Ī�L&�vtx�b� ��t�D�/��́P|�G\��J�l:\9��>��߫��BJ򗩊_hƋ�����zf�<�P~�5x9��I&�`�#`W.x��,��8?��l�A����լ�p�;-j����u�6i�&n*��O�lL���m'o�)r�L�� �Mc���t�=�=[�t���M�'� �H�ڻ]�ˉ�������֕��$�h_����Ҩ��e�tF1,xc"�E#wH��B͵���i��3	�$�!w�+� ��
;5����o@�S���7㷼�͆G�w�%}y'��ۻr�@�^|��c�k�`���f>���餜����pP�Vvgs�
F������}�V��~�]�p��Z��X�2��/�e�uZT���q39��l�� #.	�'Źԟ>O��?�����hu��)�d��W��������z:\�nͲ�E�x�I$p�dWy��ŀ7�:���]���ng�B�o���=g��^�|Z������=�+7	Ġ���-���IH�����݌��ȓ���ӫ�e�
h5���I�ze�b�u�t����;�����ga��Y�H�����\�*�I�)��_�J�&}U�U=Z���IA���� ��q)"%��5�t��a5t�z���0�F$C��|8����Sy�-�o��*~�A� Ì���N�0t����E���~�Rė/C"�;�8�m�<�-5�vi��y�}��+U�K��3��a\�FkS>����~uA�`���˗��Xw�t��Uw��/���{Q�C�5\�k��Z�+g���&��O=������e1z!s���/������r��S��S��yk�l~ߌ���d��v�-�l��0���,;4��u�O�r{����h۳q
]Gw�����`F�V#/%�4_��!䜢���E&���dݦ�C;As�]$}wtt\�~��}�լ�:P�oϨ����U�y'���w��&�b ��.�1K	r|mQ��
������|�÷!����޾B$}�D�@k[��Н[̞�K�����*9��l��q�n�N�n�iL9�W��˅D���p���C�6�3�Y�OMg��t���5^�|7\\�AO��ݻW�-��jˉ5��_�.���f������u��,����w�x�*�̷fQ&J&K����J��	1�O��WO{s�pn�g����Iߔ5^��M���y:44������m|��c�u&'��Y:�A_����aV�x���i�����ȏ�#�*�m���wOVF��Fۖ����L���;���y;3�+,:�]�5���a����gO"����R��S�\�K��*^ tv"/7�\TL��J� Z�AR*����?n��D�teGU��ג�@�[�P*#�����5�Զ��ȓK��-yj�C�K�J(��	}�����B�����g&��q�NTWx_���pi[$3/���H�̩]WJ�u��?3��Z7��`�Q��3�EPy�x=s;����l���Ձ]J�Y/٩.���K��a�����]!�F
G}(��X���H��7��ţ�GM�VT�|s��ן?c��@�<#n�'������79��=�[I�LLLnCR�>-Ss.�����M�:p-YqH�Q`��v
�8�b�c�]�JMA�&�쒗��ҮO����p�V{G�b��-[����}��9|b~��#�r22���>p�U����H_�@����MW=�z��,�hZ�kr�+��n\��u�O�8��T*�MV��j?�� �+��)��*vsf����r扬hW����-ggix�s탉B9#�{�i��o|��1���-��LS0d��S� ��|��M���)>>~�g1٨�3�:�E�i>�E?=N�x��?4f�͈��㋓�9lV�G�5�P�~��3���E���_��v����šai���1�1}���P��>ע�-}�4w���R}���L�o��(/�S�����|�~�&����3TS �7Z6�@��()*�m��Oݽrѯ���ԣ�����C&�Ĭ_��*�����/�yzz�N�4C/�7�;b]���^_���l�B>qo��;m���De�w:pv?�Ӣ��[b)�y�oHz?��J���=/�V�W�:ǰıv���5Ԗ�C��a"]���Oވ��Q���{�W����w�fR����xs������b3#I�S˹��r	��F��Y�N��j���h�������gB��eGrֈD722Z,@��~�d�jt*���͑LVB��3�b�Ƃ�;�V��� �;�>���)[�;)�XL��o�Ee힡=��[a�V]�%���|��� /���,(��a���_󅃓�J�S>}�+m/����π��k�G_�e6��:�;}>���F��j��s���G)GYi��N#&6
>��{�<"8Į����15���>Y�WTW�%tQ����﴿oM2�-G}�_�Ʃ)��a:ݯL�%2�k{�7����8�����E����dQXg�K�W05��[c�w���S�^��91z">�/j��}��c}�*�������h\/�����>�i�.C��[f�P٩=��?�Jk
�	z]|r!�^I5.W���Z�k�=xBӱy���Ƃ����'R�������>��\��*piJ=,��1qL�o>͈d\�59�G���/SG��p���E�����RT��-��Ȯ��h�?毠h�<��eA��@f��#�����H��%ޢ&8ufo�ay=���%R� HJ��֧�"1���s�(Z�Ow�m�;�{���c)�>N�EGb�?*M�U����1�������+�sWxcb�&������	sƿ��:�m�V&rؐ(��vi��%G�����*�_���¯��&��Cg�>t5�D�R��;;/Cyeg���|�y��S[I3��}�7�Jک!Q�$�X�d�yi{�-�t�M$���+8�!�8�͎N���9��(&��<�k>��,'/oι��*�������䳝����:~Tj�q���<�cv�(2,QϚ�4�5X��M�wJ$Q���M�ԟ1av	'w0l97�æ��Q�~:S����M�+kn���ʧ�R��.���݀�C������ː݉9���0������B�w�[��c���N�_�I~�G'+�l��\��x�r�Ʋ��q�7��{���v�'<�bD��Au;-d�X�n�����7hv	��|_�DI��!F�*�m���T�g9�Q��/�fH ���\Ԩ�m��?����)�-�RW��(���fF}��%ٮH.�&ek�,rg�Of�Nwб�����m��}xC�gH��CR�i��:Y�f,�#�g�'m9��}�^�^P?�=�y*A0K?�5uys`N��
+����jj�0*~���z�Qޓ/�S5np%�ŋ�wJc���q��΁��:��.�ɭ���ԓ��I��!��n��'��ɯ����e�#�?�hs�M�i	����i|�����7o�ddd����@��u(Kڡ�Evj��Ǻ��m
��v��U���tΑs~h/h!�R�:S:5���;�q(����yn�J)Q������s>D��h��X⏬p~2ğg~�|�Ľ��:��i�||x[GGJ4v��d�|u�'���W�1o��xo���FS��ʬ�,�Ƶ���Ԓؓ7����n~���#���i���R=>�z�q���ki�H�������&��boRu�t�+�Ή�&�Y�{e?�m�*P��e����g�T�-�͛�X�L�G �%�;��4�U��].ڙ��YqyiQUs����ii���R��#AKa�X�m`M�$��럾�1<�l���~�ț��Ҁ�@�侕�G����Bl)�]�����-ڋEńɲMؽ:���n0J������S�7��z�%بp�GO�۵�+�%n�?Lic_t�Y��N�$�'l&72�.WǾ�N��K����zdK98b��7�M����t:A1ث�����'��]���B���#��v�W�p��ˇ���t���5Je's쵼���Uu)�\���!�S�D�i� ;O���$��7^T�j�4g���ϼ_��>C��30�6U7D�˾K[��Ȧ�i���1��*�6^��#���4L-���kl=J%�9�  �4>�Hr�R����_���H����Ew���~��	���O������w!:'��"���L�,���U��ɒ��K �$_W�?A�5A�Y�#W�(����$�S<��M�XT�� *���5�.�8�r,�$�p���(�K^9����WA~++Z2��B���tG�+ڻ�9ө��锫#aW����PS/UZ.�,�h���V������OU���Ay�	�P�m�&D��=%�uuw/E�Wt.[�d;,Z��b��9D�y�������V�=T�m�ŋ�[q0\(iJ*y��D���P�E�f��8_���b�vb#kv�v
�xbfױɭ�j�����B��NY��,�$ߠ�^{�]���	�U}�(���>���C^^ L��x��{M�%��ɑJ3��e%���������x}Z���0�O����d�Sbs�DJ_تʮ<YZJ�@I�ݚ�A���^�L�R�M����E~H�W�
�V4���=�	�I���jI��6�_N�_�=M�'�+��:���̣X	U�����
[ZZ��)���½����� ���
���p��Š�d
��r��u`+�M�-YDGM��[TI��ꢷ�0��{�h	+E�/��3�%&&������Dl�K�4�7�q~��̓%� x��P��4�Ou�b�.�
��R���G�<����cK�=�.\�&�>&@ƴ��e�c�za���U۸��aZ��p�@KFu\�vB���3_�׸�ǹ���^���_"����RN ����·���$Z'yˁ4a�����1޶�C�mBgp9�^������p��҄�p�'��+�/_&�X=I�Eos�t�v�%��
Um*
�𱾾�<N�w�ce�ؙ,�}n:����3꾙���P����>��\�U�-��o/ٽ��[q�a�!��<iQKj���#ݽ�G=XLt9%x��$5�ϭ�e��Mid���B������p�,��Q�2y�.Z���K�;!�傴�s�v�=��t\\�J"L��BVJ��N<6�꧀�ɲ�DP�
OTvqy���U�.�?g����7��fCm	��Y	���O��+S������2xD�w���Ic�=��_�\8,���԰Sk��.N�u`��5�[f��,o��Ud�f�Z��I	� �g�2ݙ��3���]�-�4�gw��u=��]k,f����&���n'�	��� s�K���8u�su�B���#����CCC4r���>0J���c9;=9n$��)X���V���hO��=2�"γ֙�޾Ђ���''��M�C� d��xkb�}�,ࠇ"�P��;��=?m�f 6r��MX�J�DlK��֭[y���{o��'ҰV��vn$�]��B#��(�6 sL�^V9��~�������f_1Ά��H�h�{T�_H���o��� �]�܀z�r�����n!���gJX��Ӛ���o)x3��B�e��E�!m�m��4ՁoC��ˊ�(+���@yE�'��ow��=<e��t����ȵ����t�+\��_<k�M`�x���c0lx4�������	`��=ǿ�����`�y��E�������e*2,|�B)��8��p��a�H�雼>����P�%a��]���J��o���ydX��RW���̍��A�����ν��F1�x7<hL	F�Rz���i�:�p��ҹ�9�pt�x�r�0rq�G�\�#,�,��۫�6��I��n/�z�C�da�;M���-�mSCF�5�N�M
���ےdj>�(/M����c�m��D2�@{�!���[��n����;��2P��T����?;��	�|�ˏ-�U�/�4q�t�S�c�ɧ9��-H��u��Ҽ���Gg�u�ۼB�đGU�<�GV���%����Q�n�By��+�,�,��
Q=���>ӕ��y@����s��^����OU��na�V�~�E�Uʖ}�T�UTL��<�Fn�`6��;hοG�|�à��.���1'`حr�~��߄X�Hĩ��n�M��z:+�7/T��6��q�a�{��#)��DU�AP6 u�.qJ0δf?f=��{EQ�2,v�un�,����������x<ӿd��!��c?&F�7�z�*,U�n`W����vѯ�}��"g7���y��,�����~�MbqQ�����F^�;m� ��������VC�F1�����xE��U{A�D�mh�t]�����V�������0�@TΡÙEX}�mY�J�cX�XA��(f�<$���{�gBdIKޠ%³Xȸ��e`����q�N#��ڎN�PWaV'�c��j�Dӯ
�3�;U�W��66@Ex������z��`��*������`H��%���uV��Ug,�:���~���!B$���e��E7��NN�F�� KX�O5��mG70�j[��4��d��A��F*�t�~�h��޳׉��|t�tl�m���^|�XL��:,fZ��\������6c
J�(�ՙ�x����d�B�ϴ��/9}��DAц�aJiQ?�㭞\�A��{�z(R��<E�ր���"���H>��u||<�����@���D�@w���ė���;:�`��DrQ>����_�����ax�"{X��t��!OW�>�%$���/�+7� ��u�sh�����2LQ ;Q.��o�th!�\�$��yE_ۍ���M'tx+���rh�z���)�M��F1�D@���6�k�f]bIAA�r:)�iT*��7P�����X�wߩ��-�|��P3T�r);u^��~SnQ8[Z�����]lq[H��<����<I��%����*Y��^AUxҗ�'�F��R҈���8��&���7�ܼ��7�%�]�:`�����b~DЅ����E�� Pp1z�[�].7�g��#�����l`���i���.)�l��<MJ���ćXg��������[�C��Y*AA����[����}�,i�Z���{�y��ԗ$L����,��h �6	�(�=|iȥ�F Ф�	�HA�~Ɍ�q��eґ�*u��~�����G���'��UB�>�;�Y	��B߄7��a�wSL����ms@�	<�<�<��-%�a����|J��(�5S��X�����hC�U���+e�z�&�=�*�8�PJ��=#EA7Ja�E�~Z�F�0	��x�����7�,�)���N�� n�<��w!���s���W��uuum�+��JΙ&sn��,b�n}I57�_�w4T[�.���C�,|���_�D�+wz�*��Ȝ��R�4:����W�X�� �/�oP����,�i3j��U�;�Uړ	/�=�+W�Jڱs?N�5Ɩ�Z�W�!��I���mD�Y%��,��f�PGL=%�P�oO$(x���m��ᑜ*���9��:��	su��)m�ſ\��i��L��5���� �,�@ �jO�xiq�+�5�;Ɛ�^�(u� ����-	�������(jh�M�C�!7�V<��I"\�r�������I}��z�v�������}d��cVA���|�(��^jb|��H���T�%D�VqeQt·4�|N_2--�N�d�-�'�$y�pF�ʞ��q�nEI)44�@�3�}�4��6|��ڟ�(�T��D橻�m,�4t�w\W��@�!(���b�\Bݣ�t�6��#�Ԕ�W�a��+�0�wa���\�1~Ok^-�}i������ݡ�O)����bE3�>����=��Tʷ�������l���#�[Щ���r�x���{���"*��+dF�}#b@�Q�'���9)GUBLtb���Γw��c�8�JP�$F%�|���PҞ^'4�;̓F�������~\��T���
����R:�?�ڤ���%>#O2,�殍�v���+O��5?�υyh	/��w�_�[�⡛����Ax���(j�@��lP�[X�;=Ĕ.J�n��P!��v9X�u��W���1dh:Ἔ�g�3�[a�u�	`]��_���4)L��3���l#��/��A�m.ɂٸ�P�ɋ��h$�m|�i�v� �Α_�8���0ZQØz��N�9��1������?�1�TX����g�B<ǌ9�Pͤy%�d:`d���C��g4F֖�]3��/;��|n4��z�׽Y~N�]�/�(9��N9a��ԪƁd\���'����kV���J��z���/�$߶�4��"�m��@w�Kt�C�5����Mt$�=�	�Q�edd,_�������6��Ww��T��y�4�� �%޺�k��ш�m�f3q�b5����0��� KЖ�ہ��=С2��GI�,�l���A�w�igl�����}�#�s�D��N��"�M��.�`=��7��x�
|'��S�^	��VF�(���L-�*��}���r$��dJ%�vz=�����b�LZR5�p.�
���E���$�}�����-��O�a�Y���i�,���gf/{.�{2��<J���������R��Q
m�o6����+rؠ���(R�a-����������|�D��nD!��4��j�|!�\y����$P4�ps�p7Z��)�weee؛Pȅ��N�>f�h��M)�vp��Xi>{?���K�^�X����>�]����'�*�o�n�\�AE���K�9�R9f��~�pbG��gj�ccc�}222;�S��R��7h�pv�W�l�`�z ��=�B��(a�:��u�����͵7	�Sk
37��&�!��0��H��۷�Y�t1J{�W!�����ڨ�D�LU_{;	�z.dv.7�ibB�hZ�͛7!����LE�:���E�J���4�[J��w�����5�pvw���4ɐ~�4�b�k���N0�jJHK�e�j�0O}���e��4t�-)���(�d�m���![���s�e��P�uj�Nk��f��A�\{fwO�����T��Ƙ� ?6�c��G<,?	�2���CA��>����]�QMG����"^��
笠n'��������s�v�kz�j�fbb�s��H}$6�h���]�w^|e*ԙF_&�x�W�?�m~R�x�e���!���)������Wmb�F+���b��a3R��=������썞���L�d�$a��M�5�H�pq�v��LvjB$���Z��+��vTVU�>ݝ��>*�f�F����G�),zZ�ѷy.����AkX)�������|�~1�]���ߜE�#�w�,El�i ��<UX�zr:c��M��=i��2�7��!�顫��6m�������3�vF�m��U��5�
������w�X�>�,��&9��t�z�Ӵ3rg����vBfM0!-��i���&����J;�ƆJ�ƅ��;`VЋ���?	ݙ��6��}G�s�F܏�U\94��Z?K}a:#W+��Pu��b�٧����F���A�	s;����XI"�J�,`+�q�PT�d#42��³�&ub¯�?O)]�a�{�Z.�C��T�{��pl�����4� ��z��/M
���~��
���|�ֻ��� �l�)��]�._�Ltwu�NTr�tr���?+a��o��KVR��bҼ�?�z)eO6���V��Z����൫���� ��&i�If��.��C����f\Ϊv�	-��,X��J��XrD��6_@�:�M4�D�/\J2=�����K�u��s����X�6
�����������@=݄�B+0P:�z�R5�pu��c)�s����ˉ��G�m��~f�Ni�v��#S��T�$�zL�6�� �U�7�dfMMM㚫����T�9��Wz�x2�)��]�����V@��%֢K� �ǀB�
���՝�K�ma�b%�}
&��s�0M朡n��| ��>}�777��V�Aq���&��Ǐ~�Y]�n�6�.����BQM��Ho�N��}	]l�@Y�]]��xY��5`N*�-�����e#�� u��A���`K����4v�K���F��*�����D��˂��g}���x��m��@ꈻ���E:�"�'a��S����$�y�8n���Bk�u��1�դg�?̫��%U�}r*��X�ø��Bu��F1!0*���3~c8c��A��=��>::����/qu��X��y:ő��O���? 09.�����<t�����gyB��G��>u����N��,�*�N���KT�g�3T-�g��������W��L&���=4D�}�.����S���0*�A�O����|Y�W��f�Y�C/s��AVEV]Q޺���-̜>)�J{�#��_'�:�uv�nnI��;�hc�����s�'����� M_Q��6G�����2�-"��S�oa�ܽ�'�xP��[]��@��9��W{��LI���&����b��3	���wї�O���۹O��ߝ�{U�R����:�sϰ �7~m�_��n�X���i&�}Qi��R����XD?���y] �g`q$������8�(�>�u��aŬ��F��+�}R��`̍�0Ѕ6O�����իG��*_T2P�S[0�� ��m����vM��g�N�ڗ�����5K�4���r�k�t���6�z ��_�JY���i�)pM���Bۑ�nV�y��e,O�������,�n#z��Dk,�.*��io��̓�'T ��Z�F\�Α�Y��}A���?��5�g�����G���>&?�/y��{I�nC_K�C���m� ��wyys�����@oqIl%Y��'�I,H�w�9V�∪�O�^����\�}���G���t�0��)(�6`o�Em��Y�f����Nx�����4D���
�!�|��F{/*�[A`��+�#
}&��o8�?Ν��܆v;�ura����j C(�1�K�$�$�UzF�7���HF�0�(5�-�%فn4fz�mR��v����C!A��m����`��+�Ϟp'�Jt��
�d�ީ��?�����6
��l��Qj~�'�'�u�>�9��i7��O~-[X|�:b���Lz����7Bm}�J[uu�#�vB�0`��ގm."<A�����E��^��S=N�ߜ�I�fY�$�h�Vb|������j�q�|D������W�&��7��C���U�xX �m���Z�R�q���ŋs���F �o��@g������͍�>\�D|̳�r�v I���/ҷ��h�V�D&��'�B��:>!��G�|��͓�<Y������$'����5p8_�<�Rˁ*Y�lr���©N����^�wd���(�^NoQ�F�$PR"�ϡ_fwk�D>���{������K2G�D�IT/��sh���4D��H9��+/�JH�����"?��Qz��K�fD�1�u��2�����ӸCLN?��{��l�-\� �UʧqvϞ���# �觷���{R�+��_*x{�D9���DnyL ��Y	�\�Л���ԁI,e"�<}�D�����3�����}�=;ru|az`2.)ieapp�=���V蔿=W7��#}��r��h��&�������m����x!���d�&i��&���L��+-��A�O�-�\d�P�-):_x�J��͗�yw,ŕ111���,��d��]/�_���l�#dfe��(���/\�7w�B�=��8(*�I�5�4v-�F�%���#�w�z�ҿ���C�SP�����Ϧ�U���hsb�az��@%��H��Q��Ѷ�"�Zn*r�-��3���n�L�?-v�
��˟��5ꩃrBF����T�����Ν���ݥ�&�w�z#���^�`��2I �n{����ϧ��3�j��Ͱċ�A��K�ɿ��"wZW���!�>�vӌ��p�힁���������뎔�9Ӗ��n��?
*"�.���Ǐ�f�<�����Sq��8X#|K۔)V|47IK�����"�������ù��I���ߊ���<��5b����}��]O�^��QefɊ�ܦ7��,��=b�.�X}�������ɅYi�٫^�r#��H���	�8�jS�!��+!��`m�ddP�mQ��v���{���%'#��ΌI�b�qJy�����׆�}�D?G��n�hf.qu+�W�3���O�<㪢���aޗI ��ɛAk��Uk�a�n��F�x�r��M����? ��,��Lꫣ �b�}rOL��5Ð�aX\oO�G߂N��"��>Y�/�P ��=޴��CZ���xkp1�D,8U=�FR_��������
k�ۯy���¶ˢ�m,^��R������b�>���cy>�얤�=�\Ǯ�r^u���!�I��<]㟐��A�^���;\B�1���rz_SS�ι�%mܾ�	t{[P���gL.�M9��{_dK9g?K��VZ�`w��T�'�,��Va3�' `���龳�Ȉ������y������2rAW��氉H�ݗ6�L�y�>�|�KDF\삤9�nZά��r�roc3� ⋳�aaa7�a�M���"���ߘ9��,��"�;�)����%-O�hmm-IK�@�~VD���$��R8��d�d���3���勝o���"������dB
 �2w�n�6�]�*��@i���_�~9�>}^B��$on�i� Ž�xqVr��+���s����a����!����W���1V/�R��P��)o��s�\IC:��΄\��9�<@���:)4㱕Q�]��i}}R��.wff��"�,8ωv\>4������,�E�i�R�_�,���f~�a@2@�!jsW�VM��C��b	Zr�ut�A���FJ���C�<��B��
�.����ǫi7�۾y9 o��� Tzc��H���Оu*�_������$f�ȩK� ���?@7��>98�Y�6"|�4���
��zn���2�}��YȰ� �f.d�Οkՠ��vy+�>�+�]l#o�F	�
axh��C�Vs�q<��S�F́�.���杌qF+:v�A�jb��4�A����-Dٴ�i$ͧ�P[�D���������g�ك�7�}���J�W��D���jލ���-vsy!9���B��mSoN�!��|�,�~l��ɋ�XEH���ȇ�牙��Q�ǋpmZr0'''����&�+U2��99����O*����m��� K�۝�o7�x;r �����6��ɽB�/8����C���-\J��S&h��(�4uww����(A�y���t�ģ	����)����u���(�"�5�����2�0�zrкw��ŒL�_(C��x�FB�PK�ܹ�Z�����5Q<���T!!!&ox���T��ȃ���s�{�Gq��l,
S���M(�m���%j�ح���Z�oC�Ȣ��'+[�q��L$T�|D� �§�f?��+�)�S�y��Oz���P��rA��g0k����#����g�t���;@�	r��p����ae�I�*��r���
F[*��\G��Oޑ�(2��~ �~?nY��X�AQՓ�����ŴJ�Ae3��\Csss?xhߐ�2Kz�Ei���H��翧������m� �7�X�n�Þ��YK ?*���#�/��.���$*1��Dn�a�	���!�Y�2Ɨ�hJ���(EZ��夰9ҹd0@���c8� �=�Ʉ_�������L ���<99� � �1�m���S3o [�ڈ��y
)w�i4�;A�����y���E���7hIjc4�����B�����u�>��4��a�7�0�Rے_ul2��
����Ͻr��O0�tv~C]��iL�9�p��d��=� |ҎCn�z����ʯ�Ku{	����3ݗ� ݟ/�XU�B�'���n��� U�p��*�]A{�@ݦ��Β�1ǏW��7,`vl1��m�a���S��������f�<�9]}}"H�KLӟ��%�AD<@��҂�e�S����/��w2�?�>q�l�hmm�U?xpV�`�lA�-�
�>��A�}[��ks��-�%�f^�"[����}|����,�d��db��5���Q�"���9�qh�h>'�����7�l��0�yW�M�8=�ʀ����%��q�prDW�%�c�"GV��n�az^�S>c$$$�c-�V4�??E�����ʊ
����J���c �����!}�⹕O�e��=��J�������P�����Ǚe=��_�~��®M�L��~�������`�}�g�!�2G��5�����{�w@�y9:RLѓ�g1�xaD̛@���M�KHH������4������;�|��ۡ|�vd�y�d\h������.�Ԫk��R<� ��A���([�+�f��0餴����w�n0}���K}��<)����)��ME�����{u~%�0�ߴߡ'�=!��e��U���N@o�A��ӷ�Y��
@z �5�M�� Pe|C7��I���D��YB�gqi��{����?K���_ ��C����?��a���0��`�sD�6���I<��F�d�"�ws�����G��>�X����0:���1�芆��6�j��;"��sc��pG�W]��:I��$����<߼LB�m6S` R 
�yϦu����N~]+��J�C4�bv�]�ߎ
��`4x_���%J�4��r��=�����z�Vj�J��"��ʕ��j7 ��=�!��R�}�'����U��y�pqӨ����4���w�0������+�� 1(en(ʙ[�� L�N����z�u1D���w2��n{��*��C�.��a� #����NrH�i,��>�`�2�P���|5�z����K��ECt%�"���9^а�Q̡�������� �"C�����`5�0�9��I��X=$H�yD뚑h�K�M����X���0@%luu����5��C�$��N��=�ʛYWEs��.<�� f3 r�h%�:"��0d�yu~���̪�_@sh��_*�B�������I�!�ܞ�ۃ�<�V����.�C�#ȗ/]Z���}���蝍�"œ3��I��!�쉾ïE�����m�0�P@1��g���<rd�=��c�p���{��+4��K�ݶ*m�'it� 7P�$z�!����L��x����Ƚ�_ׇD���Wٰ*� aZ�O�VeC��˪&0���Z!9��[J�i]]�\`V`V��iG�z�U�ly'S��>�G��I�(��L~Q�^BQ��K.�r�:���B�����M."k�XzK�'-}�b<5t�{��vUt��d~r[�V#mo�_uQV�AJ�bs� �n� ����9HEY�����m�>7��I��.�X��~r��b�������C�9q=g�Tx�n�[�������W瘚!�$Bڜ=���o�B�R�`!� t��s!��Ͻ �΀��2�'�h	�F�Ɓ�MK�âEi��>ri�i�i��3�J.�y��t,M---E2��8�/ �'����xe�Q�z~�.<�
3J��b��P�4l7��jʊ���_��g�o�v��\}kNT\
�JeT{�rM���/m*�TY�o��s� ��@C�P����bt�5��|LXE�
s�e��o90�&��!�H�.�/�\Ho!Ĝ���J��d�rP�467g�;%W���&�Z�X�b�2߼�{g�^�N8��激��[~�NLL6�;�~��Om�'��0�}�^X1˾�p{CQ�Un����m�D����/��?����}}=������6E�Z�@���*@����8�u����TQE!SȈ�O��Ulz*��͍Oo�ܽi]?>@]��]3RD_��pォ)�=V�����pߗ���)W��gmh�Ԩ]u�1wU{�.��T�J�"�P��N�"�Ko)#��(�.~l`��� � %(F$��j�(���h��ס���������9����d�O*�8�D��O��Q	�c�{�����lyPܨ�oU��[�^�Ԭ,27��,��<�w��.Y�dRhb��(u��"6ɻ�%�\��@���K3 �Z��R��SN��q�+�{$'�.k�
�\^�{y����	���:޷�	H�e�rL;��D��3z���N�����x�6�< ß>�6,n�p�ܞ���3288H�%���;Y���I1��r9d�Cz��}�:p~�\Ԓ�5,��
�Ld�	�0%�R��a���9����R_PN{��_0F��U�U�	�jܗ�&|��z�pܳ8��P/u��_��� <Odj�����'%$�5� ���kU�șq{�&���ͱ)��7\�}�p��I� �h���k���P���? �0�U�����}�re�Fa�[�����Ew��Ukp��y�:��0ԯ=3����	�*c;PY@��&d/b�P�/�*/Z@{�?m�Gϟi�;p^ ����0�7����_���-r�k>��Y�u�Kj�Փ��+@�~����C��WZZV�1٘)���G���谂�b<FCbՋ�fEI���C�:�� JM��	�'���w��ע	oG7�K8 &R��*-Q/������1��A�dNI��A`n�o�I����"�.�G��Q���b&�l�=NM?��������>7�:�Z�����l���.rB�[��Cb�P#���#�؎�w�$Ԑ]�J&y��B�ʔo[�u���2�_�+	�W�����~�CcH"��}
/[F�����3ZW̲hT���c��!	L������Χ�8����R�����t�ӎ;v��1�RD?� �r�Sl�����8��x�9�����tP�M�>B���� ����I̒��5���8�[F��`Β�S ;�ZUy�������r�D�ߩ����:)�NxE]�8�ɃB��ݟD����-�����<f��
�ʚ
�#��&�e�8��#�?=q����&���4H�'m4�)Ed�O�gNG	�>%��ٿ@D����Iּ����Q��d<����v�c���E�c���i���ifY?f�C���9XE6�o�R2�Ѩn�M;��s����Y��� )0���=#��9�ʓ�pcS�h-<HgY_o�FU/�A�4�u��i ��w�O�@�5Q<I�vy��0C�2�H���<�g�XL���ܚ<��p��$��m��t�d��u�6��3(&�]�̑	w����Y����b&_��Peؗ�=�Jo��)--�y�����H�Ul�vh�3;��:`��N�|�g�r*g��T��
Ӿ���L* �8'J�O�8[�B�E��
0�� ���N�P!m����
���W"?��D�0�H5)2���@��f�q��О|�nG�D��������$>ޗa��C�\�b�ъ)��0����~�_dmd���D{��cR��^=�D����#�&�����p�[��Ź�� ?�B�`П�����lϣ����]h3@p# ,�sss�����jS��*p
��v�H�ʂ�S�{J������$�Bg�	��1'g�I�3Ψ�%�78�˖�����f."���A8Zan~�z��z��z��Ja0��m�X��џ��^#���}�%�3�Dw���6	���+��m�=Q�q!�(#�S1�}����>>��d��7��l.}>�諸�њ�&�d6V_!�;�P(Scِ��mݐT�4S3�������t��d�B�܈�#�c~�f瀀 "����@���>3���/-*�z���w�_��۳�c:��mr ��)!�lV�����W���F_%$Y��D-��/���t�gE(������{�7�j���ї��������x����)&�U�����1L?|���Q�Q#�2}��ɞ�UvcO��	���{���Ԃ�{Ԣ�����(]���O9Z��=�ɻ ���W�?�ȉ������6�v�ax>i��Z)xQ���0�,없u��G���|J#�:ט�c:�|�ͦ"Uc���ۨ��}���ڙaSy;m�K"3��|@�0/S�.Ϯ��Y������<�V�뗻�f��	L�0�M������L'OG���I\�B!�VFB��a��@ʛ�f㯎�'�߿_�6��x�x�5�&/OX_ut�?�yXSW�6�>�ѶZ1N`E�`�8�d��`�BFdF� �<���jD�(ATh�Id�bEP�� �2
bd����ɉ�~���w��{�?��pv�^ý���>�lQ�i��$��~�a�H�H�r�j�N��$�9,$�D���ɾř����w׬F+o��G�����[3���4{��{�:v`s�Q$z�������f��#m3��I���Źs(J��KJvμ5��;:�����{�!�
�=�I����M�՚���x��Q����m��h��hkp���a���n �peP?�Z���sYYY�.m;?��T��q��b�����;7�����ώ���vF[�8�����:��$���U�
r�9dM����EF�������{�J��/�r�}s:&6��ь��qX�3r��uK_�h�������5=9Z>L8��Ȭ�cT�Dw2����h��������ӗ�]��ëK������;�����6�L}���mY���v������S�no���ǟ�M2L�An�&
���D��dXv�Pk��б��.-��uK�;���ۓ��[6�Q�qͿ��59��a�"xpNN~zT8	~�)�i��U��>CCL'!��G']'���>F�H������/b��}�	��e�͞�7n,M�i�!���j�	(���:��>X.Y<3��a�Q$��R衼������5:�h�ɥ�w�����9��]{�z"���CC��?�ŋ�#e���n��_� �I��X''��߲*ͷ��M�4�����������zFڡbt��-��ԸH���vf�?r��DRg�_O�k�g�#K��	�5Z��_�6�VuY��]n��w�{]��Gl�EEER)���xzg����5q<`�U�SN��4�dt�;����ӟ��6]+7�
��w�\[� �<�xxF��ٻu�ɓ'��#I��L	щ���!~ꭂ�\;/95T�����O~���37�X�"��4吴�����������"���m�K�������OY�����{/�Ժ�^g?*v��p�xy{��Mpy��7gd#����]�hv.,k(�gӹ��Ш�wlP�������'b�R�A���z,�-mw�1�A�{tt��q��=vd��JIh����X^����Hc��c&�T>�5��tS�鳛�|�'�Z� �����\�G�%4لϤ�!���@�{�����8��;�Ҭ�bC�R�$�����-���m�Z(Zy�<^�% 83~�AG���˹�Qf���_|?��l5^a�� }�oJ,��M�$r �7Z}�;9m9��7]�mX6R���9�b&s�a�o�%PQh5y�[�g�H�UG�&�%�C�k|@Q�P��}�j�������};/o��\���^��rG�g��z���(�9"#�V���Z�Mo�y��<���J�m��I��+��2h�h.��f'<�O�>o/�\J�m�D�I�?W�?Z�R��ۺ��U�!�A�./�K{%B�9��æ��(��BÊ� ��_��c&��v>�-��S�jQ�~z��uѕg�`��7`�������Ѳ%�D�� ]�t5�<��L �Ti�2̵ٍ32[��<�#������$�oqm�'�ϫ�Ҫ�P��bmH͕k8�R�S������]�頻��hY�h���ݔ�h�4��"E��q���Z���4/M��`ck� �ޅ���+w��-���L�9���Pv����?��"��뫆jk�e�k�~�GHww��//6D�%Llv*��ah���T	R��� �2%�������!���Y��[e.��^��|
nG9ѿ�H�_�B��N�-B����JhKS���gF�"�ۗH���ۺ5��z�����(�N=����l�x���䌄,hBY��c�":����j���ڮR�d��u�Qc�?�Єb����c?i]���ѹ�����s�g\���Pդ���9 8WS�9��'T���EE)x�?M��z(w�8�edݒ�HT_��4�A��b�n�����,�Ԗ�R���2 ?�+6$X�!`�C���@Q�:���!���w�(��� ���bQE��S�Uo�����.��u�w�A�/��;�F��62ԼLLb�UI�=j>��>Jrrȝ*�F(��j떟�b�y�4Լ��uQ��1o��5J2x��=��Z���J�-Gx1����L7k��k�������D!R]*�9���T�}��C�^�z�<��5ڻC!mbr��PT+��&���\�j��W��n�dZ�v���ˢ��~�(�E�n/)��yad�*���O.i��GC�TԆ��4�Ri�66wՅZ�,���u��=��ak�6Q���@�//��x�Sߜ���*v+��l���ބ�U�W�r�y2>�����/؂ |�?R��a�O6T*�^{VZ�c@s}����j�,�e�)�SPL��������y�L���E
豐�L ޑ\��[e���l�s(uV��=�Ǯ�,]�D�_��PTO�O�����Fw�B��(�
J���Bd�&����P�B9[[ۛ���A�N' 8X�İJՕU�[G����1�r��6��� ��JPX�j�VDC���@�B�9DX�I&''"w�6K�;wN�Mk���2RT�K�p ���䴹��^ͯE��/_�loȰ41v}��A.�&��$-A��:�읃��ӊw��6M���qAY_6P�O���$l��[#���ޕ���,���}|r����uW�=�yEɶ'ߥNl�8�w��Z�w�3��4=o�_����d�o2ɾ5"�e�a��j�g'�&�wn�l~2�>d΍م#=��#,���l$�ܚ�V�Ҡ�U�� c=�N[�p�Q;;���_`�H�:�MQ|��FG;��+�����L���쌹zu1BO�Ug���m�L�:�3H��Ϡ`��_~izzzl���0�:N]R6x��W^Z�U�����2��<�����Qs�w�����Q�|P�q�{�lJJ��P�l����ڊే��;+���w�����؄�| �=��,|�4A�mv8��~��{4��~�j�R���nn?�>s&a]���7��^��D2D����_0���"����7�L��H��B�s�Zą��9P��'���:���J ej=�q���ڳ+U�8'�������㯡ms��,h>�=6#/oEee����t�t��� ��;Y�����	�)����ޘ����ϟ߮;xJ��H���ciAAAFF5ǩ9���J��g����ʃ�"s�Mq�*pt�CCCȈ�N��W�7b2��+�0����X�9E(G��Oc���X&Ky ���� 7��ۗ�0���A��P�����/P� ���5���D�yc���p櫰j��y�P�)@�]�����A)���T
%�.��447�CU^�b��_�j�-��a=��Z&��
����a�4��sؖ�=0�
i�~Nc�m�
33��:c�GP��s_�j�	1$���������ROf���L�vV\V��3��,ok���b,|�~�h0ǅ����ٖ��j�=�H#*:���w��TKZ��>CU*6"�m��2 #��WSm���jpj�k��� ��&�m����^�EO��˄�1�o�y�ˏeeeG]\�Bo��3L�x�@�����PM���:8;���U�˹�G�BQgQV�lls�ȏ"w͝�񿔶:���}}e	�����B�Ag'v��.4e�%A��V%An�/�� �'&%������B
_q=w���>t�6'On;+�=��wGf����?�t��`����|��/�����f��c���3Щ���w�?�JQ�����oٲ�����Q���~MY-g�p�
�S4;�P2`�S���������>/���%%��Q|���n�"�svV��
��
ԅ�#7 �S�Y5zcc���_<��h��!���d.;s挫��"��B�+#����XQc~��֊p��������h�u�sԽ7��}l�ԍp�546�C��
Z�E�LmEQ\��.������R&��i�� ��+W�B�K��C轍��4
��eF�g\=O�w�ȅ��)��^�q(M��CyCP67���!,��{�"˜�U�6�=�G��]�_�����@X�:4��!6`��Wv���54���'��d�fdli���>�|�9�1#'G266�j�����q�q�"����z�C�r�޾+o蜤bY{�Q��k���i����=������#(���Z&!���|��ڈ�2�J ��xj�ʕ+�����]S�TJ������.\� %-��x%i�v 0����G5gfFK���Eb�ő<0�����I
$�/G�� ^[vɒ%[���P�<S�����ii���$CD	(��e�z
>������i�p����88l<}��Qk�c)SrPWI�Z���2�2����i����K�Z�9��ޖ�u�9%ӎh�*�]x4 @ыe��IT���ǐѡÕ��уy��wzM%���99��2x�5x����"��e�%��*��+��F�x+pY�`�%A���������ֶ��ు#���{F&�	�&��I�?}�P,_�rM]vժpD�P��Q P2.�}�d�UH<�DoDDԍz	�Y�cЮ�x{�v�0��-	��NP���B1���%3��I���nY4/D��[�PB�c`@	K���C��P��"N�-~H1.�+Fz&+͋Ԗ/_�ޔ玲���<�s��i���)���wRS'��ii�tx_�b�����s,c��*�j��x���[�n]���Q����ɧ#���{	�Z��`�rd"�Rh�j���u����|����!Zr����_=��s�2��			��R�ԉ����@4LfѢ�`�%�^*�X�W�J�[����yn?����om���)'��bhz�
Z�1��O�b+O�I��j�h��I�i�B*A�EC#`1��D������zFn�v�4k��g��x8�<���x����zFo�Q���uy������ݻ�'N���׷9~|`�S����Le�0�PD N��X*�A��-��1�Wo �@��E/w��M"���K���

������	���~E�|�_}AQ���!�kc1n�(vxG���d�[W�jkˢ�J�٭����<Ӕ�&�uz�nގ>f�����`���_�A@N���e��**o��P��\K�$mG@f��Z�������1m�O����ً��j�]�^�&��q[��K�-�Qύ�=��Fb���&��ޫ@���+{�����F��1әj���rI!��ޔ�1�������-}�wo�B�=iZ��Wz>?i��]u���T{p��cG(��,SD��z�� zN�`���%p�P�B����a�Yש1�x��o�*c���dZh;C����MN�l�ܹ��nZ.�Mٸw��3c� �y��}���f��+��q`2G�ׅ�$�����>����p����
�������!V�_�xQ�_Z2#��>���1��eY-}4O���YV��u��8�*�n��3��b�^6;�,��XҸ�}u�����L���$����3�OK�q������Z�	SN�Kj��͌:X!�]?���r�-�B��,�<w3fS��{+o�;&�z���P�K��d�;kr��S-�̭�{h�\�K�vKz�Wʡɒ�kb-�nh-�ܹs��ڛT���x�%�D ����k�\��bQ�Eu��ES���:f�৫�����n����#�[��M`��m3���Q��VP#��ɼ����f����8�\ӑH�����@���n��!`b���������4���ETg�R�x�<�{��F�v�?�2�h�U�۸{]���t�����/�t<��,�^3�Y�7�0^���x�k�FV)u'���}ҳE��mv� ���{@Z�t���:��4%�X����Co�@/��B�{,z3f�{���L�NF���>�&��m��]�Zp�������AE�c�����$�x�4�����<�kXE��·C̺}�^�RhnԩK�'uܕ�����l���3��?��(Ċ	�f��u5�	��)��]�:�b������
�&hU���,٘��<�Ӆ~'���b��xF�&���"�fb"�ewo�i���on��'k-[��?.Z.��1�>�:�����q`i�!;v�N}�!����k �86����~{����̺��r*����Afݎ�u���EW�\)Ki!�l|���!J�˜�q���~�;$Kzf2Ug˧��\7׈>�:��^S*����M��j�w��JX��� Y���ؘ��ð?����+�$(���v(��g�+B��z�����_.~���○_.~���○�]�l��<�p_.~�����&ǂ?�ƿ
�W��X!�|xQ�W�/��|���˧/��|���˧/��|���˧/��|���˧/��|���SHCސB�`����ݹz��&��w>^��|�-��Wت��N�Ν�=j�V��),�n)��9�t����[�Q�ϩ]_��8,����_5^��=f�M·֡?�^�ݓ�7�v^��r{���oߢ�?Gӄ�����(�{��z�T���/���R�������������I��'� � U�`ݶ�������~�杰�q3���Ʒ�j��g.�Ő���l[��қ�|��!��C]]y�=<F��7�B����B��/�吪*-��"�������$� %i��6������|��-�I��4G��-=�Iڈ�
wʙ{����.O�r:h��9>M� R,�v7Au!���?�e�#𦯵�翺yY�u����?ۺ˫@Qd�σ3tBΘ�>�����_��i{9�&�9�r�5�\^�Q;Z�h��[��:�">��*��C�^R&!+�f@}�E�9B��ϒ����I4�������?��������:�
݁�E����'Hy]Z�uNQ"HqK�O��W����"%�u�h.k>y�Mj�x���;����3;�7���M��`��{��k�T��!��- ��uujτ/!�C�XdZ�<~�vH�=kw	|��E[|��/��Z<�R����b�H�tCbӝ}��1SwA^?���g�l�ӄ�gE���t�]K���N��ލ�ݻW{�*4�_�������~�������^x5��a��b���K�#��FdL3j����N|�w�p��0���z沃������m��y�{M��~b��9�*El]�g v�	|�׊����\O~�.1��S�ߩ	��|��*M�b�M�ޞ]�0#���g1���?44$q۶���z�q�֭[�%`Q��V��
���G���bQ�
�ñg����1RNJJJZ-ŏp�K����!c�I�8%�ڮ��������Еb�|!��^'ш���>48�c����9$���v�Fm����J��w@S|��������鯲����	FEPq1�3(��7e�`M_�6���}�����}�}���>�z�����LjP��hA����2��{Q`��SRS���K7p���job%^Y*��Ou��Q;����o��W/�W�z���c���G�R��Əa�6]A
]��@���+��Ж'� �d6_b�B��8��%��8v옾���(D���]�Y�`36�M��MॶLd��+��wy=+@֖��������sZ%�.��Q���Y�����?�< kS&�!A1sI��7?����mXPI�~&�N�6���_"�'���W��%d�$b�Ow�2�ד�َV�q�*=��p48*������~s� B�["8Z[LL�X�P�����T�kE�I�XZ��K�]��v,P�i�Xd���jv�M_�M._.)��X�^�2#�4h�#.9��z�*�e�_��0��/��E��i}�T���^#�:�ho�X��o��Q|�l�+,�z�C2�WQ����h�~T�q���®��~�:���]��,�M�{/���e;��,�w>|�LصClW��`�0�"96��S_UD�� N�ӂ������Z!�j8 #d��-��8���?�ˏ?ϼ2w�+Ne�֡��TH��h�`�Ka�cc�5�� ^�6y���嫒�nv�B���<wx��Ŭ��\�������-v�;�z���d�.YH6璂a�&�E$�+��w����rW�q�L��ܷ����h�u��2,,��F�Ɠ�s"���k���֑f�M�Y�#1�~�Yݿ�aI�y��n��z����Qm���7�8��p�ޝ
���!z�$�˖&t8!ҡ�v�BJȷَ�g	�m�F{X�
�������m$���ߞw��7~JJ�$�����V2�uw8C��lֻ8&��b���"��CNt���.fu��YU[{�<��������s{웝F��x�ʑAud:�]�(�:�����s9�S�A��%�1x+��ա�x���'�O��u���Ѻ�+:��.\�c�Ĉ�����K�E�:���"���M�w8	�K����L����#�1BH^FC�`��fvcoK.��3B�ޣ"�$���C��������I�C��t���zp�������zSzvI������!GHQ��*����ڔͰlV��%r��*Q����j̠�#�L�r�e*�1O�1OԢ�5�a�U{d���D�\pNd��C��H�+N��9�Yw����"u��	CJ�ur�ѫ�n��B���.{�'����l�(�V���G�p8J��L����c��dait�v]��?ڧ��� >Ml?y��l����v���-�و>�	�NK���Q3f�>b�C�r�`)м6��1=���	��;����K	o���n#}��ź�:m:m��v8;4z�kK�����%}��>��e':6/�������`�DO�B����-L�R8H��k�86D6�jұQK���<)�� ��n�e��M��^�J�������O~�z�c�Q%h܀��W�S�=C�*ۻ��߈>�	�:�&Կ�Ʀ����w�L����V(�L���̞w'bR�%����]0�ӧO7E[x�J�i�.��}ߜ��[��!�߂c���D�s�%���7u��i����(i�ouy��x�X.(����ˣ5�/;�J&���ry���l�qn"��`���5�'�㝰#��Jƻu~s���{_��z�Y�e�LD9Si����Lv�
���W�%��aH֐$�_\}NCz���߰&������հF���N�@��YE��ty$�ꋲK��
�_Z�����nXD�8���M�t S�}��F/5���i<t���*��Y�?L&�6:F)�|�� ؼ��(�� .�t�K 9剚���Oq&��#��"i0�cD�B	,�%*�~s(^6�����6A�)��m��s�<��	Y�����:���)����q�����v �x:m$��$����6�1��<�A'�_�|��ZK~��i�v��R�\UB4�kI������ۍ	��{Ж��9���gn�sA]��-Mٽ�7	����No^�-0�qƏI�KZ�F��
�ۇ�ޢ��Ĳ۳/O��;�&͝i}��S��3駺k��/�*(�<4���P�Zɹy3L��+���0�޺mυ��9����|��,Nյ��3���i�0����4�Y����w�%M�u�1*R�0�0��Ǣ�޽{���!�$Ϝ��@-��nt��I��؊�FJB<¿�h4�ƭC�5N�k.H������	�������b%��ܸrc&�&�q24��� �
s!9fC�s��*��j;4��i��@�����ʊ\���9*�Y
qt��F��%	CJ���N-]���,YB�S��r&��5���ڗ/_jeܿ?����}2���i��I0��������$���4B�yA[��w��p���':ke�\�޼~�>��.��MB��� ű��w3��R+"j�/�{31���{@ӓ��
\3y%��	}�w��j��h'W��+��PN>z�H�`�-"~���?q�]�����w�z��j�"�d��znTpc�8Z��;��L��+�$;cL��ǯAk���H,I6lG�i�C"&�PW�����]	ۯAF��_wx'�q� ���d��j�B�)�eA�h�tZ�d38��Qq#۱�n���4�i���N2�]�Z�}��'�y<A��C8�0=�.�嫞�Ç���Kn�p��F�Q�6?A������Jr����v�~���@��l%n�TE��Ũ�G$�=(�v�CMM�/� |k�E�}|wӻz�L�gR�S�EV${��1�Nл��r~��K�����_ze��ݗi�,dƍ��l�k�	�ȝ����)��i�?@h��4Ӹ��'y�v��MM��ٙ��S�d	h����c���i]���j�ˉ�������A^NɢԘmD���(���D��EZ����>�����X��8�*�ᑀ��ޕ�[i��\v,���`~�~���.����/Bͅ�cmE�QK��Zl��`r�[��5��g?61*��Ba�Yl� 2��<6�ei_g����V˸~d��H���}drz�;�e���G;��&!�<R�{P�y��<��.ȼ��p���N��{Z�d��R�D�(��z�ѻ�f;��poL��G�+���Aiw��Uvo D�R��2&��!L�S[ѓ��p���J*��ǜyZ����urZ]�n!Z̏�d~!�}3�ۊ6���P�-nVb�H��^�`P���FR������ׯW���!�$"��Y+Jۮ��z�����Bi?�=�3}hk٨c��UG;�1�7�2����C��i,�K�» !��!Ӹ�l��&�V�&���T�"����nU�֊rɾ8'�/���9�p�I�yML�삤�tٍ����X\��]y���C� .//��[8���3�Z �4F�DY�29�˨@��R���~�/�v��B$r�Fj％�c{�]{�5���!��0�ג��Mh�&�D���3SLk� ���F�7�3��P�W������8y;O�������n''m62��Ԟh��=�)�Iu�cED���꯳�
��c	��IS������,�U����f|�v�l�;�XG'r>���F�VT-��Y�Cm�J+`����x�G���Zx��x�Q�AsFz�@���H�}��˞,�Xkd6��D���y�E���*�ԑ�'j���J����&��hn�BJX�.�	0RO��M*���uE�i��P�g�:le=r�u�#�ni'g(�1;ژ�Y�~f	bE×�V455=a����N:�Xi���Y�=��pʐPft0333s,���v")�v��iUU�>�r��.[=~amz��tAἁ��Fe��3
Q�F����Y}�t��3�qsP|���k߲֝����c9��}�iWd�qW܋��>ZDV�g�쪯e�k~B;�+�c���d^V	����G;�ʙY��		_��W���Y`d��M��T��T�����*KX�Q��w�3=m�;���.�޼iS�$��Q��mȝg����p�B���r�8��t�A�I�.[(�1��.�GFp�1�3F�o�o��y�����WL[_<V��ڳ�CJu'ù�8-��"�I���p**&�PP�[@Z݈�d�� ��o�?N�z����{�ky�w\����'jV���L.�xد�=�32S�/d���!�#�]�챀�~�ظߡ��"��!#$���%��g�<������hoIl���������+�&�;tZ`aj�&�*}9��N�N��	Z����	Ov�1�I��7^�k�
�Wډ�h�z�wb���n'�˝��^�tZ\�-�^_%����+��r�$����%�����(����v��/�Z��!X����	�r�Q'�*����ۈ,K��_b���d�]����F����lR?R����1e��7]Y��:4�ot��co%|s����<
C��$��܂ſm��������|������B�8����,徖:�煝����������ӃA�p������D�S|�;�D|eψdapSk��I�ȝ:���:M���c��]qP�����	A(�⸲i�@(��s��L�;���ߦ#2D�zڻD'��M��ˮ�y`��{c�Wճ��z�
���(2%S��Jl{g�kE��O��E�+:<��aKC��U��0�l0y�`��y��p�Dfuͽ���s$O�Z��)}�Ԟ:择�\���i�KǇo��0�hTDB}ϴ��9V�������IE��AD�!K�g�j�@�£�r��$�!����cI�|�#NP.�����~��,^)W���̠%r[�[ᔾyx&x�\�Fx-Ӌ�g"�B�ĊZg��v��/<5O��RT����
g��)؋���N��V��0m3L�?����9��:�k����J��~�t��r3w!@w~%�e��x�]1*H<��bv��9��~�o�����q�1N�] �2ΐ�^p�ҟ%����Uuj(�B�DCI:���wF�=��}ѽ�V�*�;_+������?~��-�D~_��_r��޶�♈ C����ُ�5k/��&#�����C��a3vװ(���އ�^�Ȳ���D����)$�y�N=�c��"��cG\k8k�X�\�&�B��K��Ђg�-��c���r��~�K��J<S�g���:Q��Rsz9C�W��SO�#�N-&`y����OD��X��U����e��C��.�)ii��u��Q�^`��<����a��dB���뙰r(�e�C��h.++C�ύ$��4K�u�L�]��vE�!�4gtr:M��]<�mC���bj�%R�s�����8Y�Z����!6����O��q.6޳<�gb:��l�V�2�Lf?�U�<+�����V�q��w碚Nʐ�6j�Xc�x�� -����;LLG�D�{U89�&g�����c�N4�VTT<$"�Rd땐˼uK{��i�s�����a,�yJ��N(��Qv��2-Ea���j�i"�2r{��T�r�RĢRf��z*�:�1�y�!2d֡)@����U�ȼ;M����\�/�
��R�F��0w�[��U<ގ��33�������*�.��bټ�5?��x}��d�!~��=����ZȐUnР�J@����CD�+6G���n�͗N9V��ޗ�1�$�Y�`�U�8�x����gW�Yb����B��QI��.��F ^7i,3�}�t�!��<-с�}[��J��S��#VM��K��2��a�ݑ#o�ހ
�'�����8��]s�ξ�76�gg���N�|��S��K�O ��o�=W�\魼H�U@���y��~y`���F]�L:l%�2V{�$K}��u���P��N�A���+-�����������i������֒�&v��tP	�@�p�M������ڣ��\v���w�<-�/G�$mO�|(u���>�ܟ��3�6�S����w7"���d��i(���/݋������kll,��ZԊ��U�S��p���T�4EU�?j�� J��ѦNv����֦��Y����WeO�i�k;����k�����(�jPI'>�v� i�gh/��w#z	��=x�,]àaH�V�]���_�������T!δ.GI��"���Lt�!�ۡ��y�9��PBKT�I�xZ�6�Ȋ�k�@���`�`���N��%�cl�����C�VrE�����Q�&9��ۼ�	v�Il���{%��q�nk%G�u�ʪu	����#Tc�\K]�h4&��_I~��/�W�ASAN��v('�����oe��~�
1뢭��e��A�H0�=�z���l.\^�� �t�%����@��� ���[2O֧��y�f���t=9�Ξ��h�RgD�1�i\�p��XȌB6�S�.)��x�tK������GԄ�sO=�/6�-��}�+K�"�ڇ��?p��k���̍ı�����?�̑2��~찑�\OUi����d|����c�S��U5�u�]0Wq��|r�,�7�~b�Lò�E�❮��港G4�TE�n���,���/4��~�Z��sӴ=�?S��V|�i�Y �?8C-($k7r��FFFVJH�\!��� �P"�Ÿ^���ר1�I��j��A'��Y�Q ����Ij��?C3���)m�F|�&q���sO%E�間���W�2���b�s��%5�UCS���1�*����}5�&����D�+�Fw(?�^"=���gտ��4F��5���ҽ�N�9��I��m�|II��2%�O�ٍ�;�޽-�Qi��Oΐ���OU��u�p����=����o�!ghH^kL�r��R�%IXp��<�����!�O�+�X�i��Z70`n��Y�66�&Z�	.B�Y�3����*h��0F������ϱ�7�|�[��6�n�4v�y��b�t����Dʡuy�2l�l�K�a�܇����`��>�G�z��k��3 *��-����wN�($�|L�y0�v|�]S����K��X|dH�a~s�j��kbX�Ӫ����C1abĸ�"�o9��_���V`W�:J,I�>�M�$���ơ,m���Lï4N$���z?L��\�X�gv������� �I�SG��H�|���(�쀪ТV9���X'�Ơ�����5挲��Au�Zr�ZR���yv�Y���[�T\v%�	��&�>�e"��ZQ����XY�(������fS��*n�.�"�Eh^*����(=MWptphҒ^���Z�y�7��^���X��CY�X��0��F�C�dp�j�@
��1�=�%�ɒ����gN9���W�c�cIL洛��	rJ���f���U��4��8|�gA�q";uR��M�}���M���{OU.��%�C����uu�q��=%��t�w	��*ӮZxf�|�V;w)5Mj�\m��s�q�d�~i��7�3��[ڊ�~u�����&�v U�E k��9b�@�}��h�����=*g�'e�=�6�4��@�����2�944�oab��Ig���I��i��z�2�b���L�SNkν{�c0����.e@s�5��$(rr�zL��h_LD���z�%�f(M�Eӝw/�c5	���ށ��ÁTW;P�;j,?��VM"o=ȭ��ق:�s�qTbELH���7y�32S��l�3eC��#J���TG�o��CC\����f��#X���m� ��%%��S{Ʊ��Ȧ�Ä�Ɇ$�����W������t�~�z��xW��%J���(�r�8��*h������ͽ�Dy�nN�t?u�q�T�&�Nk�"�P�����!�1377W��a��������}v]]]9f��H�0��G��VV��:M`����u����#4�8���)��3ќ!o�RY��m2��iP#�ac����N�u;��Y%��krVR�����9Tr��;�n�\#�vYd	�X�&�����d��-�H��p(�!�6	|�k��M�4��-���``���D�(۽�"A(�wi����ɳ��<�J=�����	���Y'S�lo��*������;��-]���Yo���Z2��M�+��Kk{FR�ъx�V�H�JN�ݻ��⭜����)�gD�|�@����"����Q�?�+��뷹\n��~����*�`d�`<����&�kG�\P��
�`#"<��yB���sqm�OE4����2�����2TY�r�Ni�B�w��o�J�?�5OFI<��s�˷�O��.���O�eT��"X�ho"��D�:��"�"f�e���L?�\�����䴨��'!qįh�|�?D[������yvc7Q��O)e��)�%�Kշ���g^�q�)A��%�$(3M���-����y�U/�yZZJJs	��XBcf���T$1Je�{d��ܘ���~6j�#(��]����������qq�°jBdI�6!�k�����qI��X�|�$�j����x���555�׎����R���=ȰV�Iy���N�_t���f�s�\���ڟ��l�7<��貖��Vԏ�	ԣw���c�6�F!W$�m����p��]�&�Wj�C���J�tel��DKօd@-q�����C���"����C���$l�b��r��[���L#X%��r9��U`�}�D����`t���(&��[ԥX2�z�CdA���	��W���)��{3�v[ٝoτ�ƃ���3D�ǜ��[����8"d��Qo_�ײ�ں���~�e_���p��8�p|����z=��[��o��}$f�pU�����Qm\��E�6`�ȠK��:�b�u�P�\��K�1G�\GnFĜ���_M(<}A*ݱ
����U��?������&օ.�By�Du����F���:o���֯�����cx�8�O� �[��P�l��C�z'�^�=QJF�D�넢 ��/���0�1�r*�S��S�����>�и������DF�-V�:F}eY�Xx�{�A���-�6:���j�j�p=��Cw�����(�5�<g�&��~�w��V��#ԟ,��n���$�K�Qȥ���{��z '%�+��zZh�d���m��h��n�Ih`��\mHp�#� ��5�O���K��ވ���,��{����r��E��	���
�!A]�H���FZ�<�o�Y�ΘQ[����y�|.��R_���t4!�Y��y��b}���ȑ7#�V��k.��[�"��r��#��%��)�kG���#bioo���^�.�:OM�7�J��DQ@�!�-j�s��%An�(1RjB��7�����$�mK�����eH�͡��lv��O��j�vF)_6˧���>TF��o�y�5�~����ˠN�;;v,���9"����[N������J�t��Ut�v��`|����N�.	�yė�B	i�'�R����̴��t���D�zW>�~�x�P(lՔZ���%!�]RF S��g�щ�ΐ�<	������H�����'��G1;]�!T���')(v��יh�*�tQ���&_��X�O{����過Y�֕2�?�;��r�djC7P5�5�(ʵ��q��?85O� �-Y��M���)�^���xH13�Ǖ�=��������؆�4nS��b8+g�o9�9�)fh#���%�[���_<��gЍ	)@�9g���)Ą� �õ��YE�갅_��Ox^ I(:
�"H�����=�ë�r퇴[��oJÏLf
�{^�^�r������<�!��Ƙ����j�JR��\1�%�~��gup7�A,b�I��K����s/V��#~�~�&p��E�#��;�i�Ԅ���#��~� �.�>��x�׽�@�y B�ie�I�����T��V��<��z9���A8�w�(6�{�ՄSOY��w%��v�=��ۼ�U�g�n��@[�?Zrܾ�"���`֩C-^+w�g�(��8�_?Frn��	�<v�tK��X:a$X=�k+&�"�����LN���Q0~Vk�/�21����5���w�ʵ+�	�7Cb�Df�Lie���'�!�Rpْ��cפ /L�5�Ί�6}��Q�u�%r���NN��萷�8¿>li9�������"�z�憦��z2��g�(kK�]�*��Y��>���H_��'�uے��#��{��S�jB��*,������c.��j��A���P�7�U��c34�_��j�Dp�u�C����@�\Ǵ���~�"THّ]�K�	G�{�����!*����)��ܽjj,�`oo�	 Zǽ��(ĨR-��»y���"�9��������i��n"�%8e�%��"%%%�qJ�o�_������P̢�~b)�9���"ەl��ty<�_i��va�[hÚ�r����~�U��������z6��y욡�˗�n�1��$� �ju� ���֒�\�.���<Ra#n�#Y#D(�I�_�N�Ԑ�N<��X�M��Rt* �ҕjVۡ�<�N���(�qC�k?K��rqee�5fG�Tr*۝��W���h ��tP�zt��x��)���32L/AA��a�[}��ک�P��@n�Q���X�8�s(y��:� ��B��goQ�đ̪d�N+�	��X����l���x�]�܏��5���@F���')>�=�����y���5�"@0�r�A� X@��i:�]�3������(��0��$�!�A�����J�3���[��~�)(&�&�6
'I�r9��<�evM��Q�����e�/_>���K����.�m��ur�U�K�S�����9�__�?\�5!�,�]�r�X�g6P���Vm�߈S�xo-��t�Vvיڍ��^�����D��jFzZ5���j8�uM
���䜈��@�1
ـQ��2��]:S�I�ѱ��ԓf��j��o"*d�\ ~r��q����j�:�s[1iH�x
>�+Q�/��ȿ��G�{(IM� �*�B6\ܻ9������V�vLN�7�������-��M�=~6�}ͳۄ�E��@����.k�*oB	�Y�,,��>�/�	�쯾3A�h� A���Dm�E'�b/g�Sܙ&=$��z�Y�,�>.j�Fn=��Ҥ\e��"�W�kį$�1��:�����)X��"tN� F��f���ꖢ ��:O��>���Z���X�r����/��^s��]��P��\�#��=�{8�i��{�$�~<�λ��7~��<d��۫O�&����e�O�G�{Q��=�u��v���U�{-��7���3��U(�9N9�v����1�"ף��	*�w��|�w�������0k�..�Y끅�!��n%��n, J"%5UKNN�ƽ4��(3'߽�ʸ����u?�u���~H�/X>���	v��N�ՒPns�'�x�;�@�AM�)�ދ 1&S��(-���,�Ă��A��k?���,��i��hg�RL�SV&�_���r��h��"v����F�y���(��i���:���rDkk`�wtoH�8����Ī���&����l�n&��~h���XD����PUy�	������ce�g��:���I��K�@�(����%�a,E̺�G-������ߠ���g��Lf���F9-Slv����yE����A��3����'�̲9Q�����Ch�_e&qZ��V�z�5��/1�����%Z�����ה�.ҍ;��>��Ri��Ҍ?ˮ1���a����>��z�@�I��T�S�+��zk�v�<yc%��3�������Q}_�mv�Rd�w�[t����5Ǩ��(��J ia�Ĭ�2�J-^�:~Q& N��i����8ik�_�֙u'�.�����5a��w��V�1�aw!{�5Hk�]1s���	�S执��?~����g4�`�L�offf�	�C�q�\�bC	�]K]n&�R\����گ�6�&IJiyw~�oyĪHCZ�M�q���:`��w�O��R<w�U�ps����V�9�������b��ݓ�ĠW�������í7.c/!$g��g�C�4���g��w�m�Lz�5W;w�;9̺D>N*$��׫u����j�X:mz,j��ɗ�a�g���Z�_v��IN�v֦\� ��_�����;��v@ʿϮ��O�d$�NNo�ѯ�B�:�s��ū�.�r�ϻGK�&�f��=(6vin{�C���f��ࣜ��M���{�7��g����������i[_�Z6(����!�5�"�E�@D�@�~�}ĉ#��3XQ@�(q4,Q�FQ��o̍>�R�7��{��{���~,���2�Ӕ����w5�j�
}��D��=�!��H��eR�R==�H�Q�/ef�?���nD����|��_Q���<��!���O����u�Ɖ"��~��:v��Α(v�U���&=��j��,\qL��)�4-qJ���`q�:z�␈��� E�
�Q	a[�l;����*\���A2�ˎ�X��N(���u6m���8��bVֈ;xZw���׏����^���θd���p7,s+�5��'%��8�U%b�8�fr33��!+�Q���[&���1���!D��K����#Ʌ�\�o��a+@[�˵�e�da�.Y	���X�ҟ�`ہ'oWh�-T���*ZNNNk��J��9����,\�Dת�(�>U�Y/r��p��4MF�=�?�|-vlԏ�U��J��!'w�J�w�Ĕc+�%��/)»8ΐ{�J  ^ 
�>F��_l;���O��:@�BZU��w��ۋ�Jm*���Օ6Μ<�t-��LƭǞɻ6�YB����X�
�c5�	>�K)�Tff��8��:��4��z���٣��@�o�lNff�K���k�\|�~���Ɓ�V4{R�MI�߸q��''����0���au�K���@�%*f��C���$��������t1�({����3����>����?�Fg#d	9��F_M2������5{y�o� o^� �ݭ{Fă�'df����V��H��Zs�\���ɠs�XK᛿x�~�w�]�C"�N]�G��-��eӣc�7�r�Y�jH�,�^�?�N�͜����!�`M��~��u����~�����Č�Bg5�3_���݇����W �����๳|w<�qi?���Gw��n&���?K�ea��ZW�L��f�k �O���+�Kܔ���sY��wtc��#�1O R�@�[G0�o��A?(��V�g���.I]t�#���[��E���L��v�&��1pk�k�z��	4��Ix�����O��V//�ALL9�
W��q�;_��U^�+M�������l������[���7�KJ�&��+|ޏ�� ���>��AV��ݹ���CD��_��v����"{ֽ�i��j�b�.z��E,��,?��
J�/���.�u�yw�\�?X��!nT�2���{�8ՃD�������D-ӐW����n��AF*�i)��lȝ�ַ�9����<<�$V:�v�JP�x�-��y���?Rec����u�_�RH�dK.Z����7�!I�H�v�����[����l[�N���]�����>���t���\�="׳�J�mҷ�޽یΠq��v�ƃ�6��c�ݤI{���Y���+�H_�u��g7��3)-���mA�J[Jcq��$Դ�k�g�����}Tԍ��Is�Q�E�^��F�e�>?בF==g9��Az2��p;�m	K�Ŗ��糥�7 �lG!���?�2��3<��`���t~����D9������l���|+��X��+�O��)`M<d��<^,�i][��	�RZ �FOP�̟|||�YWH���n�D�5JT��[!Wc��s�&v�%���gpLS__�J�]
������NG�$� �A�S�b�����u����nz�+j����Z��!�~Q(�|-�`�f�6�7�����~xH-�[Q䠦��چ]q��85[$*�I*@<d7��9#����(1����v�$0��DY��[�f6�p�b!��1��� G�M?/{�RÌ�I�Q�)���H��2���N:R���|��e�&q��n���?y�~}Bqa�Ǐn����z^~8G7B���.h��R�uFo;���f0�;"%�}H��:���E�*�����,f$F��U��7��
�u��@����%�N��O�+:21o2M;��7E�����n��n�g�u��r����v����y8��k���4������C��ʬ�&:�[�"��� y:��>� {�b"��n�]nۑ?3.$O�L�~Ȕ�O��xU^Y�c�G9��ƭ$��6���[�-�7���p��9x �U���
�������]���� "�&w�o�<$�`ڜ�����y�Ђh������
��Syi�K
&R'���Č��G+��L�m&c�-+�|�6���̧�F.=���1`���JP��¦�>I�V�av����&�����o	�U�ڎ�R��_�~��<=�@E4&C��i��p��a�j�u�y/����|>��v����iW� �𫦙�d]]4g1�k�Q�ێ���x���4���t,�~�Dq�F�t#�g���%5l�F�-��ִɊ��;T
�����Eާv^��7�x�+4r�P˔��h݅ǑCX�Dt�i$ܘ�Y�����;��j���;�<���J��1ߙ�25�7��hX�����Q�ω,�c��5��|>���G�:��{Ď�Es!�cSe�O�(�d<�]q��{䄋����.���%K�78>n7�61��qW������u���B��3 :��Ш!o�k^�ΦBfے��q�.d�3�M�M�!���ˤ!��I�L�ސ�~XM[�m2W�2�ʳ�	�O�>�F���I��b#`�
H�W����i�*�ã`��8��3].���M�9���MͰ���
��^��a���{x���.:E�;��%�P3�\l���0�I��m�1z��v��jժA�kw�r>C`p�'Y��d�|I<�������D�L��
�ƀ`0�Fz�Zm�I�+v�)����F�O`��YO�2����t5F>j�F=�P�2���(|��?Ě���6\ugG�ye�i���ш��=��"$�a6����� ��5���oY����#`�|޻p�,�oH�0J�VyG�C��sS{<x��(|�P�]:�;��b[[}6o~v%a��IW�q����O���������酹i!M�bz��L�������۰�g8m���]����
�5z�B��%��H�0����A6B���A �Y��k��r�,^=����Si��◔��q�#c1_joAmU3�'������33[V�ܾc$����)���lm�S��[�m�2g1�Qc'Ǽ��44���D���uq[R�c����Sxu�X��b�e���m@u,�m�����t�a�:�DY2�'p}��Qt.�`��J�l$5����� �;<ǅ���L�&<E�p���).���]1����FF��l��E�Y��v�4���f{���GqNGtR'·Z�`yH�-�s?r�X5�h+o*�	
���5xֺ����&���&3i��?Rv���/�����f*J�Tr$�p�E<$���au�v�t�^D�9�3�q�� �e��[�ϔ[uE~�<��(%����3&f�2�}�mSp�v��w�ܙ���9�ʁ�~E<���kܓe"���^$������^[Ϧ"g+9!�_�Z���e�12��`���z��`����6��Tf��0��A�`��P�1S����mY�z�]�$ FNsS��UHa���f�X�:���j����r4���utԫ1s`_���n5l+X|�j/q��߄���2uȣL�͚�F��0����l������q�]�a�b���&P�'~��E[�wq��	�T`��uUl���ׯ��%���R�D@�ϵ��ۖ�Ӏ�1�7&������F�m�
xS��� 8��V���y�zL$��S�0<��I�Fb�33��Uj��1Te4�(�vj�"���+3��c?�J6��W��Axq��H�Wf��Ԅ��]�.ŝ[��_�-��= ���\M%�kyE�Ak�K�������.���������&��:؝�?Lh)i�;U.�}��Y�����'�n�[�D�rO¤��6���.q��vu2.�-(��H��(��=�g�ʹ@��l���� ��L�tt�6f�'�,�~�p}5b��JJ�����tTB�[=g����Ss���Xﺉ�F�b1�`-	�uu�3���2�Z���|6b��� �=��b^�*&�N��B��<�ሒ7#˵���?�%V��ӳ<��T>l�Z|� Hј�e���kF��(em��8v5/�k͎����(y6
�3#v��D
��^͎�#j�yYYY��P�䐑R��s��
S�Ջ�U�7��[М#YmhO��gΌ�c��e� ���:�NDyY��˦MÅ�ù�\\���m��- 7mA�H�4����Yr�y���K������s
D-f��K��6	C1(5��׮�KblFn�n01�|��(%9je�6�������^%!5����X���D�+�����,ᾤ?���`>K�0�m,�s]T�K8'f��\�tZ�H���Bz�%��[�ʶA�n�c"r�< ��D�%6B��`��S��؂5��E����n�^��~�SQ�5(����ŦBC�?#��s��G�����Tnʗ�J���pu����#[�(4��Ex�]��j�D8�>³�lL�+���"�h�D����|�B�������D�X��P�������9a���n|We�F�da��+��AXm������@��_J���=1��]�[?�g��^���� �}�����.�5��=��y�n���"5ݲ/S!��}��m��kD ��}���DL�D���CeuU���kK���;����19ݥ8�@�-�˒�,�aFM�lCi�s^J��Ơ�{xk������O��<�������~4���.�DY(`s���s�Cm;1ziE{��en  v�-WZ�TZcrB�1-��`\9'��hJ������OR<�ƚ9窐����*Y�pb�E�^�z{�J�궉�u�B�9�,�_��\�}^�q�m#eo�$z�>	6PԷN�@ّ�괤��H��j�:�e�J�$X�)h�E0�8ÒF��u��Q��qZKs�xQ壝��5�WC(/OO�4F66��?{�v���N�nlf�a���1�p�4�X��ȇx����$��ppuՌ�z��H0bl�>�Q�),J���ˏ���'�Ho5Y��Bf���`[���z�mG:��D|�َRݏ0��c� �P�>�*�CL�
㊅�$]^a���t�����()��i?�iN�-��c����?~r�.E�K��� `� �$�ϟE��vA!r�2�l������j��e���^�N�M�kE��ҕ��T�YIW78�'��s]����?�-�;mؐ���E�8O[��>�b��7!�o�ݾV��յps4�cmŞ��H�ZQ5��� |!��[�;
��![�c��6PU~�8��u
�U��S��3�Wc�����x9ZZa���k��������e�����8�ۈ9�o��9��h�Y؇��uA��ӯ\�rvس�Ѹ;㳒�Z������~��ne�"f���þa/�œ�*Fg���N�e��:���;G+�����vV��ʟ~�G&8�=���z+Ȟjh�
�m`P�&ƫ��ܧZ\�{B����X�H���s��I��A2��qS�_�ό>Y�'@;S�ѝ�Gh<0�����T�8a�'ħ^�6J,�c�wx���v��n_'h���K�(�O}���aQ����;��ow@��B�D�b�q�+��P�G�޽����E��UbZ������4�z�  �^ 73�3�#�ع�7|x����F�i�`�zM3ng�eБQ�w9�CbdZ�q����~���~I��PΓ��m1��u9g�5���	��R�B�<ؑ�����H�h7��u�w~E�<�� !���$Ƌ����4���l!��jo��GSccT,{x���)O�PV�$����q��}�p�o��nᎧ�!Ğuqv����Z�����s������+�g��f��ƺ�k3w�R�� .5F�������{�"��nK��d�C���5��ëن��Twf�AᑶQ���X�Wz�Z��w�T��`*o������!�#�p`�q@��7B|����ŋ����X��6��T�Ǉ�ʅ�==�/��I�����	R]d5�~�s�S��*G�,մt��Ml,���]��Rn�i���x޻� �@��(xO�$��xC��?�
��+N>����d�F����lݹ�i,fz5�\���_���DBD�f�]����L��|)''�	�JyS	���C�B�
��|a���O&�4�a$�}��^�IQ'����J��͑�b`��GR�>�
wU����wt��p�X���4v��e5Ht��*?II��7�̶?Pz]���ll"�
h
�1oY lTg�"���95ƹ�<`�@�^;kv��^W�M\��A�3n2z�Q$�?�O�*Z�SF��7��4�֕�Sl�8���_�mt�MCv�~��{m��G4?�}�e�O��opPݤ�C�O�e顇��#�Wv��?��昋��	�_�1QD祪��?���dD�fj��t�~8����|��n��q�>���u��ٔ
L!���AGky�QY�ME�e �����砞�k}��0W{�-��XJ>�n:�<�=�p���O�QB � P��d�\��q ��F�J#[�E��P�y���%ާldz1B�.v,�_T鈎�^ɫ�������ZЋd/!�-%D�����T���;+w��&�Ֆ5�D���έ��Q���0��>�v�Þ楩$ܔ0۞�"N�֜(1E �1�ˇ}}}�A>����0T�,�!�@�v�?6��.�N��%*$�2�
���{�2�@V�;�&|�tP�h5�/k�����Բ,�D��N�z3&��������Y�������B���]$�Ի8�@8�\Z�6Q�>.��ZʴH9����Z醡�� 3z����Ӳ�aT�n��ea�..�,���=d�x�߇�_6�#��y�N�����%�5�`4�����1�j��K�=��;7�B6>^�7U����y]q�8��܆�BP��ۻC��3�!�_-@}2�$�ڥ3���&�ɖwJ5WV����7�c=��K}F�j���o�}[�D�w��7� [�r�n��/B���F���d��f���p8�����= 3�σ�o@�	d�#��Y�%�3���7\��O���u�Oָ���^mn�h���YVh/�_�
T122��ɷ��A�f��{�ғ~��m?Y�����Z��+�I,�U=K$��ϴ@c7h�B6}2�&�q;���>��w�קԓ�XZA�f�ɪ��U�ވ�#�"y%8���ぎ���l;���켼<�j��&1�`�2�oh˫��^�k\�Gf	��0h���#o��vY�u�l��3h����U�����V-`��<�_�~��e/�n7g�[�A�\��í�?�]����Y�A���i�?(q����a�d���֭�Gy�4��ڞW%�"�;D��]!�;�Ʈ؎s[E�s���婜e�Rͱe��QdJ<�����ib�f�L6��P"@����b�a���]�3'OP�� ��G�h�c�t���Q�����q&$�R��`ڌ^;�^���&ʕ�@���S<��u!��?���|5��<���5p)�?K&IT���Av�$����o�H�4%�f<�S�[��9ΚU���@����7{�K�^�Q���}��LZ���^���r$��|v�����i�j���4�s��s~��4<�[��^�7��L�>o�(CUC���9:������0\/%;��Ejj� ���0X����>>>swf�!����կxx/�3�;���P2�zHi��Z^�܌f������˗��ə�A�gO�xդ�m�~L�� gr�4�t;x\K[֠X�s�2 �:900���; 37��v�$�9���S�6�վh��+����� ���ՠ7�������2u�-�ϴ�8��a������\�ja���0�_ET��s�%Kzy���<r����R�UM�{�Ǧ�9U\�Z���D(=��q��w��/��I��!y��#�)������Wo���Uq���٢_9��?PK   .��Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   �z�X�ة� � /   images/8e621aff-3cab-4d84-92e8-90ee5aaf6d75.png4Zct]]�Mnl'76۶��F�ƶm�qc�qc�N�_�o���>?�^{,̵�<gG*+J!������!�H��~�a``���_OF �̯�EUJ�f���LF\D����/�������zje ��} �,"
^K�v6:
6�q3:* �6�@|P��FED8a�K�AM鵷y
6�9�k�q˓��s4.�����{b�7�sR�������r�xm����	5���x=�$	VI��\Ҳ��L��6E����ZܘTIy�c��4n����bO�������'z�<�Q�w�ڹ�[�@��p���UܧJd��ʑ�T&���Ϝ�F�\�|��Q�Ώ�o��������M���NIg~�5-K�??�-����;��C�Y ʥ�W�8����xڋ��G�K)��Sq�U:	RBt�O���eP.��rΧ��3��nN�~�]�%���L����9g9~�@�a��z�Z,�'���[��"@�aW(5!��X���d����z�-3�c6�,��T������P+�);�0Bg��|a1�_`�@~���b����'�D<M��V 9����-��\��:�	Јh
Y�P�}��d��ƭ�;n�+[�Y�{��9�y8���Z�������^��lG�k�I���o�]W[N!p�]/�Ur>���I���,	� ��9v��/�^;)F� 1���u3�UT�_���#����������ڟ\��ܫ�8����͑�v�����{Mw�	�ם�㳹�qu�c�)`e��/6:Q���/zɮ���� L�p�<���,ב��v���G���ڹ!��G�'q����Z%Y��1�]��ޕ�r?�)��t-&��]�5���� r@��h�y)v�;�?r`�D46��U?�F��?"��hʧɲ�gl����bŲ������O� _� �ƣ�n�1�5��T�<���u����d�Bm��JGq5tj��Xl>�}3s ���ےB��<5O�e���HS�y?�>�-nw�n�2�S��~R�q���k��k�$	UT���n|�{;��5;�y��Ñg�
����,r�vc�ߠ�Cvχ��1�����ٸ=@Iĝ��Pb�.&a	ݫ�&���|��|�����6���P ��i����u04R��pM;��.*d"�T���b[�4Be�\`�G>���z��̓�����y~�:�h�Ϋ̅*�-��􄒈�S�u�Ɛ Ih[T�U%�w�+�'{~5p�?|��wv��Y��*�y�8���5�p�j�k��&x�i1�I'!"�C#��Q+M}�/�
Լ��js����a#3�]�+*i�4c%���
dLɱ�ط���[��Ϲ�QQ�z	��+w?�w�xyt-�if��ǆ�	�&CM2�Y�D�Z@�:�k+Z�F`�=�Y��Ώ��]�,�ޘj:,T.DVy���7���!AE=��u�D�&;���A������c����H�6L�T����f������}&�5:|��5��FF.����7z"c#�Q�vvfQ�}����W�g�"��q+�ϲ���[c������$.#��x��ސ���S6�jA�Qx	�@�rG"��R��{���S�U���x`���x���[�R��N�Qw�\�5Z�L�h>4
���/�%�x�7V�u� �,˝SFe���Å��� ���v���!|�-.�oE���?9]Պse� �\��찾�db�`̢|�M�A$�s�?O�	�gw���%�y��u�ʵ�s�ړ�1G/�f��?�q߮�#�OР����2�حg3V�!��`ȳ����tr*I+Hǰ��s�M��̮K�;8;f��:��u?��j^�q�F���'N-".���Z�o�`]|���s�Ƀ�F҄a�I�67��6d*�0
���r���5zT1�c&��~�B!O����L�`9h�SV�9'�T�<~��R��TEEERο)%ï�,
�������j�����j6���z�-lgK"�ڢ�"��n0��MV*�e�~/��yX\&����[���f��fQLLLL�Mr� mM� M��U�|����#O��8���~�E���{,ZbF�v���J�a��h9��6� )���v�X�b��w�!L�u?���Jn>]"��;���2���b�N�"����\#��w�:�M��?S��?�ɿl5��|�����.����cL��?b���D�E������E<�:��r{���,��H���50��^�XMC�����d�	�_#�����A���6a8r�Q��o�;ڒ�������l�ۆZ֖:p5^ȯ�\����Q8�az�0�+�c{m4��[æg�|W��JYx�M_�.�j����s .�h5XK{��&��!�A��l�{P�Q�'@D���ڟ�y��ّ��|������q��n�d���c���#����i��0�9ԅM��n�-NI:�d$I���ta��̽���$6�<F����@Ny&�=�D���f�������z\��'@�&�Bl�c�RC)�h�����;t4T��]�1 ��6�4 
���P%&5:�L�%x�٩}�UUltD�+]�&�9�7��	I��e���*g��kb�4�'�=N-_1�/�Iqt���)��B�7/[�T�/���N�����ҭ����or�u;�Hs��p1	���&��t[k���F���G?�K���Mi;u(2[<�zg�T+c���*�4�z���J���*TԶ_��Y���^��=��D��1@����NMK
V���]S���,u&��qÅ�^�4��m?M�5�չ����&�|��O�>@�r�����72��]k��y�#�����+�W���&.�O�����,C�8o�D��Y*A�ê>t�Y8G��^�B���N�Iؿ+pq*���Dw���2��aH�hhp��9�ξQE�����>�|B��>����>���[�ya�����;84�lM����$����J%}��$-
+Ga!_��@wI^��IVlF�$"W8�Q$�I�}��pJw�M!��?�YU]a�/������W_8��苙���ҰP�N�6/z�he�������(�*�%�"Nv��R�����@�&��݄��Q�Y}��.ܗIʌ0��}�����W�x����#o���X0-�>����F�~��;�8"P<KV�)�"I4E7	�
��+4�r �M���TBr5�g͎���U����Q�Y&�g�-�:�3�9���K�^�4,p"��*6�J2[�0��e""-�!&^�\��6�� �eb��r�Y@�\��l��C���}a5"�Z�ʎaE@�KL��M �������F�t2�:�pA{����pRI0�$�h$�Y �Kd�K쥮�������DI��AQN�T�v���ɜ�R��׀H�M��/�PW�זv��D�]�Ѱ��,�+���I��T��u�):��de=�h�H��}�(���qK�h�!���w)��Io�C����s#���q+l���$	�~@�0�r�nt��{O��6�S�L�^���"��<�Vj�����F���<|�^ry��p����|��P�0;�1��*6�]��Nl`���Ѐ2ҝ���L��'.��B���oo0�dk��l���+p��m��d|	�ߢ���n��-/����=����?���W�����O���!cn��1��~�nڰ[M�@ 6�<\l��U�~�ol�D-��cZ-?e(ANaŒ8G���w^nmK,?֨����z^/��V����.`���VZmǦ�Ă�k-�d��g"�uڄ�������jLH���� �<�|^W�~R���V|�H��+��)�8,L߫v����t�*�o90h���M�G�/nޣX�7�;'��n�{D�n���F����9�A���ōy�n剌������o��]���3�O]+S׺�U5����}��G���2·�n�н6�`F�o��4m6K�l�
U��	��!~����%C��L�@I0��ﴸ@�-4���l�WO�b�����>#�p1	l�7�T�aH߆Au��}0�	W�-���N��%SB]l��6].g�}o��j�+���5-�s���^,��,�"K��{ c,�Nb��[�y���+4��~���h��Ԋv���#[��D����21$�n����8c�5�Q�ѥ������Ui�U��]�����g��3�` ��bEt�u��I����鶱����j��r�뽲��l�]|ɸ�8��4&]�s��:����_���/�yT�;��x9��!�0ZK��b���/�'�pEma�܁�E���y��Q���4)�����'��`�S<!_K�r�iz��G#��d�j[�������XG�p��l��e��|-�.�a�>��4�Ð�vޝ��_�o�������f�z۲�	��@���J��Zˏ�ƛ-�S}����\O�)�^��ndM�&��&믺��� ���.`�nz2t=�+�E��e��n��[{=.���5�wd�3�K�������»�4H�ۮ�X���1�:5t. �Ǡ�ş�m5Lgԟ1��`Iк�����p>���x� ����G�����^���d3��zI� �)���x��*g(Ģ�� ��"��&k������􆾶2u;et_r���8�D{7Ϸtl|(6���0CU��$�X��qfj��B,Ds���{<�I|a���\(&���4�=�j&�֗^6b����v3��u=�o���#���]d�1�������e8�Fa _���/I�wO��8�S�ߺ��?�_�Ϫ�l��Y�à@�_�m�K?�y8��yd�}��`ID���*�ϗg����n���B�jΙ�bD�����Z��R���)�k�*4 ʹ�>Ë� �$�S�4���tCL�5���y�S���ƺʌ/ �db���j��u[:�#��{���������s�q�[��b����R�3���܍����" �	��{)8�bp����
nr���������l*�*�h��`�;~�nX��o�f*�����AI��Q����.�i9?���oK��7�O
�Lh$���/;��q������:���>����zpF8��=�xC��{���uu0p6�|JIIa]�S��9S��X����r����,�H�Eҭ��0���Y�=� ���`���B��82�����7��	�|n���{kT<�N��3��l�PŻc��'��p�Dd�7%P�,G��~o�/����7�t��C$��:i�K�;<��
s����cw��26�h�ӵ�ï^e�l�Q��)����xG%����^
׫+9��A����8X>РA��7��R��8�������1��䴖���B�7k�]�Ͷ�-Xc��V�`W����/\r���z.{�_jGC|1^0��y�����9�eD��${!�Kat?���׹PB��0Vz�����t3���LB�s6R����;���o�?$��[��T�h�������E�ea���L�����p�\*.ǉ#�a��VM*�34@d���
GE3�H�&�mk�G�sL1�M}���8��"��G@0������C�Rʋ�n�_轤���~x�s�a1^gꭾ�^9���f�U̅���K���D�L�ewI9�k�;�e.�~���9^��#t�]��0ŷ^�
��������K�/L�455m��K���2��ٽ�����>�"i�<��nd�A�r�p���YXƕ��z�N���:���TR������V�o�H��|����D!<��Т �p�}�	����M�4�^����V�>�ߟnl�����w���+��5	�FD<֫���ȗZ�˵2�/������7�,ty����������� �ǐ4�d������Xu��ٖcBFΦ4�p��W�d=�+��={�����R_a���[g,���L��Mжo��(�6&�#JƼ]����i���b���_��-������@a�"��r$՛�Q}Ѱ������V��/>"dڶ6V����f��d��`csZY�ŶrA��5����yt����&�!��c�N|*�)#E�~6Q-�2DI���ݛ��j5b܂��H�.��q�1gLR���0�;/���ɀL���"�?,c�W�|� j��b�%o���W<��?�:.q��=n�~�� c*�r�D�q,�_�u�V8UֿX!*�؄;�7������U!��l:r[`�V�C�l�o�)\�K)��0�v�wi�y��	�Yv�]�}y���i@��d*:�ʐI͕.sb�#�h���%X�B՘�O�Ӝ��:�����G�)�|1,'�U�8�����N��:Z�$�����*N�A�i�C���*�gZb���C���@4���

�}f"��<��]��{���ֵF_AC=�H��ߚ�*z��(���[m�m�C���������9��d|��}��v��`bη]�L8j�s?��uy������ר��Ld�3�X���|N}���ÝLw�������p��siA@4��{�g�H��M׵�,l.�N��Ơ��[�7]��=)Sʯ��D�]�J5z=#E���b9��r����<%fZ)dF`��d�Z�C{��{�m/�p7�H)y��N �uW:��1֞@)�٥��z�"�����7��\�_�3l��w��"t��dG��ZK|(R�N��%%!9r%PA����-��������6�к��h���E����]UV�o>2Af,��p���."#`h����l���"�y��@S��*j��<��e�)�8��&Ȕ/R�{���jCmOG����?
�II{_ܜk&(�k*������`jh�iXG���l,��M�w�$�O���o��ttx��u>'8�M�����~�/��[y�6��v�E���&��t�f�����9F/����Z��{kD�~�f�JJ%��!��f	��=U���q����Xr@=���+�9��\�U�Lq�٨/h�+�G�~S��%��$�����.~U���X��,�)Q��$��UV��5��[f���쮐�-Z)�d�I���P��M���r;s���lv:��F��9,V�j�ֻ��]�������{Nl�D7e��{=_�F�y�3Z��޺�2Ԯ��X�9%�xT�մ9��tj��vE�$��~�wBq�\,6�5x�a8+bw��y�*�_��<M�� �X,'s$���;N=$�A`�W!鯁md� W}k!�g���ʑ�U�
�eC5+.R�8����T�'��ð��5��}h~V[x&`�:�i��>��e	x?���~챹��3r�O�"i2���`d'ʈ�^^��������a�1���f�[������n�OV�lۇ�0$|�p���T��/<'͑�2�w���Onfi���[w�سJZcG^
�#��>^B��z��'^K5����לG�RB���;#��21���/I���j��F
�y��|_�������s'�k�{�6 �Q��Y(�H(`����,LZ��4��J�1��?����s�^Y�+=��G���D��m�у�Q�Z`N:�R�5[��	zaT��+T�2G�S�� X�E�#�8���Y*�J�ac�
����8���G�a|����y~��K���T%h�#Ho{�ER�|�w��bL/��������9��h�(f��%� ��	��9Ŗ?�������6�?��-s�L2�E��f�	>�r��1�p��A�� ���	�j��ʼ�Ȼd��p�>��\��ǈ^�\}e�A���g/��/��~~���f���]a�=�-���	�1�87�x��p�a�E��~F4q� ����+C��_���#/�3qD�ԁH^��L�C��s��>���.{O�}�[9mJ�/��f�z'��떬�.aR�eh�AOD��by��αyp��(��
�S���u����_���'�2]\����l�*�>o���{�B&�z�b�ΜeBn�{�l�o����+���#~N�р�9�7�Oq��#�cLK��`Ez�U
H���'�"y�JcddtT��{�4t����0���Ip�"��O�_�'S)Z	�=uf1D��.�+���)�r����
	w�G*����*g�T�tw��x\T�rG	�Q(6�$�m�
�|zeT�����C!����`_�0��pN$��"�@>O�>��T��屼���T̘e�~���&����袂횰�Swn� �����K{y�n�%tlK�U��n8�����u�^�<>�-0{�!�!Nn��+�{m�g�S&U���k'|�����m�!��\1:g�LC�I�����5��
O�X�w4�F7�Z�]�C�|�[�� >jp	��,�Ң��Dh>ѿy|�@�k_:�F�Oy/�^?����8]��><C�oA=?nQ�����}	j"4������z��>7�
�ys�Q�+�I{w�������n~��z�3�}�L���M!t��h.1�?��������ƿ�n�������]�p��X���W�H=����u��2U��<��u�3L��ks4V0���+���Ԛ�'��f����۴T���h<��[e�}�������p����Ȥ��6>W��C^��ԑ�^�`�p�Ç��c�,"�U����ް�С}�XчըT��B�s�;`������=�c��ӧ��zi'�0"h9f�;��{�L�6]�U�����}Œ����?������F�<���Q(�F_ߎ �
�o(�<��-�>[aXV=�34�p���BFͣ!��Rs�\o����Z��z��zR�q3�}˿[;�[��)�����k0�M�l҇A�����{����t�o��g�jH�����N�m�[xN\��f�-�_�w�]��A�WN*u���L�e��Ó�r"O�9�[K��y?�k�FjK!�g�ѿ}��-5Ԧ�_�p@�����ݭ�t}���!3�ϼvk��B�8��F������Gb����U�a���w�����رR��},��'8�{��P5#�ft���5�:9¾��x� ��x��P�\q�����"Z6��F�;�R��n���{0�57�$�Ӟr�+��4Ň�y��`�d4��� �D�4�L"jz�H\dus�߼�P�<
�c����D�6�=����<t�D�a��L*���x�2W_����J}u�Ο	kab����4b�R�{�����z�!���`�}�K���ߜ+�3qR��UmE����H�EZ@OӞOe󀽚�R�e{�0"2�ze��*�K"4�j��x��|����,��5x�8C��"�����Qnu�]���h&6�U��m�
<^�vn�U��6�Q5��������	�f����	}al#��QM����f����M�)-�&j�B<�P�=�,���G;{#��:�HO�;��"ϯ�=���Ѡ:����Cϙ��ُFaI�)��t��Ym�qj~<���{�ӽ��y3���B�p�mk�G%z.5����!=$$,b�-d��e�����,�G�?=����I*�*`�*�*����J� mUs�.�@��x.���63;7$
z��*^�)��65��Nl:�j��a��m��rPJ;�svɆ@�9��U#�C��X���ڢ�m�������zG�+(���G� :4zM/Z�q[�i�W(ɡ"�ߙa�B����g6ח���C���H���b,��X���$�:��~�`���)[0���}�IA�H�{�d�27�VyybYp�°�_K#G��9	X�4�n�b��vgj=�EAMy#![�~�ZV��HJ%	H�"���.FMHv��;=e'Nő@o�x4�"JI��Y[E����Rp�z�E��(���J���]��H��T�l��NC�ҊZ�}��o�U��t�j`�k���s/��1Nd{O"��弧�J�y���޾�>*�W0�n��Y[re:8J�i���Kۻ1nI�׫�v�S]��uR��Іղ������[[/��OEU��ʰ[�FƧ"�D��P���*s�D[��B�l���}	g8��&E��� F߬�S���} �9�U¤F�����d��"D6:.���	0]�<|q�NZW�8�:���@�Ӑ �>kҶ�I�!s�o�8�^E�}��T��V��N>D����l��%�%��\�SP�(��y"P����u��d �g�+��o��(��|��A��WV�ڰ᷃�H�#1�q�$*/�"&��߾��d�>� ex�w�+jm�V������h�s���S��Cb��"��aA�v�,�ʒ�&�Q�f�K�Z���r���eW,{[,�&� �L��tkts���u2�H�l��'a^"���O�e$bh�y��z����#�r���%v�����J�sLFC� �+�|��98(?H���u�\B.�����N���+1I��_��&��A�6R�K�ʨ}`i����d���N�"D�uL�2��023�Z�a�h���=�B�iF��������� �fy����l>�ro7����h�:O��}{���>�q,v'��F�t��p�������,Y:�!c��Yga�tM�~6Y{ڌdF��j?�������z`֒�s�n`�5j.G�"�G���@>�Ó��KF:�J��u�f4���ϡ�F�>�]�v���Š�8�#� u���\��჉��q_r,bD&�v&7��.6�� B���.�e�N���g�'�<� �;O��%�qL��⟞t�-9��=�+X�n��pI�'��"1+�!��RS �oy�	�k�ޝ�ߝFs)�f
x;eo�QWw��Bq����C�!��^d|��b�*6�T���]◦T�KG�\`A�_�d[������,*�ތ)��-̒f��n�n��$�L#T�,�H{CK�O�- �P5�iE`�ᬾ
�TP��O�������n���G�(��
qIǱ��H�wC��_�;ϐE�4		�;[�9�˝'���+[��x����Xf�D���y�5�Tc�GrX��a�d�ϑ1>�z8����#�rH����М=|�̦ˇ_���� ��9Jħټ~?�Ġq��3D�-�өfbp�}�A���:P��i�=�v��\	~\�����p7���b$:��d�[箷 �%ʐ�ܮ��3]0�K����H�ĕ}{��Ps�P�Kn��2?df1�3����шT��
Z��w|3L!�X u�7���x��e�EN��T��9�Ŵ����AH:		�Ce�F{�������;�<�A��J�v�Y�\���n�|�+�׺�}	�.!�̇ëἳ��.E0��$A���'�_Pa�2ܭg��?>�
�й�i�ڻY�X�42��&}3�VDZ11�h

K,�8�CE������~5�`:n�o�$Cdj�-���3�	�!���Ա�/�C�z�z(`�d8��(Ig%���@jm�U�a<�;�0` 3�Ϡ5>QT˷n�a#h�S'� �Y�(�I���xKF�ЪX.u��*����̤@$��+(�K� ܵ�:��S�f0��!��t��p&�\���8���-��[hB�^�n���dC�(�\M3��l�FX�\3 ,5���*�2�;Nj,���p�ߑ���?��}�;�缀�f��,&�"��5 �M<l[�pΣ���Xب����E5����u��GΝ$YL��6��@���W�ʍ���s$5��NP�eޏ�ȅ��Q���Ytϟ �HN���o�>'��<�i:���d��?u4�`u���ko#) Ϝ��ʨw�n��´	��������#����CB�ӳ$BpH��uPW�0<h��t"��­�����,ǒ=��Q'�Ht��ۀ
J %,pY´t	����p�0#L��x��3�c��g\�|U�V�	lV��)�WD���L}<��0��#FƟj�R%�e&XmH%��U~�����s��kk�p7�ª�B���7䂄���A��T7;��HO �$K�<�*��d az�=d��چ;�E@�Re��܄�ǺbE�`%%�s�Cf�;�- d�
��a��<��G�3��;	B�4�-D���	��j�rE�V��wY�������ѯWZ ��6$`��h!�K���y�,�*�#�F�q�Cf}��4����b����V�E���x�X��nH,!�#�{u���{:�`���������4G�*���ī�w(��*��=�Я/� 2,�Q�͞<ee���}��sX�|��/S�3˵{�#{S����N=k������� "X��@���M��UNB�f���&��F8r�"�a���N�x�1P�aR�٬�qY:PX�X�(�]��vZ4%�Рz�����1��#�Ư-�C�]a���L�1xa�Q�W6`n"9	�� {�r�p�l$7����C�'�n0�TH��JG|�c2Oj���2š���FG_#�����\�K���^����|�҄�7@��}��=V�|>���fnm�2S� ]uY S���=�9E�+W��mr,��M��r_)^$V�
:�ˁZ���+Aݓ��G���w'l�5�N��NG�Q$���(N�[g��Nҍ�����+H�+լ���t�rzh�7�7]�+�Hٚp�p�*;��9�Ɖ������Y�qG}N��`�heq�������vŭH��@�(!�[���N��U����Tf~1n��#��
���v*�~���kb?�n�#aC�MPh�i��ō��k%o�Σ�/ꂄ�FW(C��@��}�I+C��~�#ubAn����}**!>T�[=I��r�+��EI1��i�c��C��5�"G����D0�`݀	�'NN�.Ͽ�FbOQ�8��$9qpb���:z^�	Y,1=TJ�s�o�����pb�� u��?�v�5�����ٞ�B�����$���X;A8�A#"|n�j/�ʯ�Q�+�u	��T��Z照E�(��^�\P\>j��F�%� �0Jى8[8���D�����m��Byh���,�4x��E������Vm��>�H�3&ռ_78\�
��]����� ��&N�i�ۖ"*��>D^a n[�<��4P����:g\�0l'��)��]�f�� �l�c7�&�X���<F�<>����DRʂ5���VhiՅ�CuZ�O:��~$&:)N�nr�:Wյ�j����M2/���'Q̙em�0O$�'z"Y !\��4 Ǭ��'\A��㑱-��`G5�RS�2����[��,׃�L�W���U*��ۓK2� �]�Y��f�Θ���u��@���kʱB��WE�&��p̐hn2!DW�K-�WZ�H�k�u ��f�����w��6��O57�F/�e��"R �+��΀�j�]�&n�H@ Thf6NP�O�X��w�w�sJ��KYe����T'�"zNA"�k,-�6v`eƉ�ȁI�pQYb@"$�Ql�<�������]XXǒ>�v�V�����	�=M��#:��j	�i��i/�r$��5��Z�{��'�к��.�u�, �����x�ca6!�0:b��Q�,�.9�Ƽ��*{��n�5r��CF4K+W!�e��:�(Vo~[���X��x�~X&�*� =�VI���p�����AQ!�uL~?Vy��ƞvX�<�no�¨D����w�ΗPN\�ه -��HE?H}�s@�]|�0���3�A��H	�qߛP���(3�qi	�b�M��M��>�;�I�:����R\*�]�����2��|��l�~e��-#֩��Tu4e���8�J�xN��mGִq1��|q@�V�>�_�-)��˞D��8���P��4��,T��Oy�i���B���N��B����/
M�z8+Hy���#я_�Δz�}m4�����F3�]�Ʋ��E�VQ8�άn�\s��s���JF{��芬529G�E�`?{�Sa��`F�D!�Ѫ�����/ i&�,�ZU�v�<��f����S=9e��K6���_���4���I���	D(�
�&�Cu�IP�X����E���OSz��@� �\�
��-�ʔ�9A8�guT�)R`�R:*�^b$7�%fD�άԼ�?�.�0�(C�hA�Ϳ`���4I����ZŨN#"Ii�e�S���\�hq���<��7K�0*��-W�|�؀�k�����j3rIڐj/cG:xO�,��`,O�\��6��YU#�¯'=x�u�G�����q(�jhSBI�hJ�2(�:�+�r�$�@���8y��r��c����^��!kR���J�	S,��d�m���]�X�mD�b���#JL<E�B2�6ȴ�+8���/�$�DMd�I�񒬼d8Dph i�~�:�1���	�H��{�Y7*V��uI?�"u�B"��4h{n�����"� ���M����Ȅ@Fki��,��L�\�N,.�2�R��K��u��S��:[i�O�a���h�x�qH�Y� k{"��C\��&�-�^؇<���_p2�-*z(�}��':aJk$Y�}ή�A9�/Ԋ=%� ��c{ W �IJ �I��-���x�8C	�h����b����0���)z!?3�LO�����Fç��ˉ$N_�M=%���TTCu�$��B8
g�N8IWi�p��X����jy�@V��'� �8�L�ʁ��Iq�i���%��q�"B�E�씹]�T#��זXf�<���;cq2�VRLp3U!�EYCj)�U���K���a�X��[�#�)�\��E3��I )8����{��^Pf�1c]=}�ݹ(8g$�U�=� �������{�̮�+<��6T9���;*wmf�����?"6,aa�dk~����e�&C
>�0��Z���o�M�y�%�H�d���V�0A-�̹#C5I8���? m���23w����[go�=u�pc���~N���y�C)���M�������6~@�&��*�_��Љ�����̿bn�hK�M   p�P��_1�s&�*tAK��;�%xJo\Ir�s��n}6<ҧ�j������H�ԲK�(��k�����R�
X*�!�^˭)��@���ɸV���A�<	Q��c��j�B��G�={4,3��<��o�TΒ���~]���ַ��������� �89^XG(���:vNbb!ºr��Z���Pn}����w��xUz	j`D�T� �XQ"��T:�Y}�_�=D���&��޻��񳼪r�4so����zweuY��'�b醙j,dn�b�l��F��|��zZ	ъ��X��94����ɘj&����C�elRZ��ct�b��}�G���[O,_�!���,����p8+�峱1F�PJ�fJ��1�������Oe ֞9�� �|`//�Ѵ�9�Z�ʶ�hGU>��m+l�h	^����9�,=�aU��3��)�6d'4{��`$�ݎ���8wX��;{o�Y^,�����?�R){�He���WB��) ˵B�{����~M�Djk����ԗ"g;jL�V�z�֑�i#���'�[������u� 0-Aɑ+Hb��� ����ѳD�WWߩ~�J��S��gNMʼ*�xh���V�$��eH�[�`����%_X<�Q���1��ǝ��e�S��
���� ã����)�)�f�/�ή<���J���UHz���LBj�$8����xT��v�өf�^W���4�%��G�f����T\�2Ѓ����۹��$�/`�w'YN1ezE��{��QJ{����𓛔��-2d��bG�!%��V��'��c���-R��.�IۧwC��J[���?�� K�8"���(�T<�}!�)ؓL�=�_������I/�� ����2pt����*1PJN	G���Z�q�ߩ�kv�m�o����v�J+5kj[�AQ*	�X�Ҁ1�b�?6E��L��)ƌ`6c��D)<@�+(F����^U����"�7mZ���M�� n=}I['�
�d���B�N��>1����z�%W˱������V��Mc}�����67r�D^j?>:����9@�v-��bf���mj��՛��g�k�����@�$���ڑ��h���^i���X�<�r*i�5��"��M�w���+���*+�Ý���)@ێ�?����ea$3]zC�}���h	������0������k��ջ��� �D}�@]
Ji�
�G�y�m��8VZZ�
v�",�r�"d�u�Bu3 ]N��B@���U��p��� s*����l�>��WQgU^}ĖB�:�v�)���.��yW0�n7�)��E�� � 5@ʿ��4v`�����2���Dp����� ��F�IƧPX[I�����x�dl�lA�,��U�(«i����A���̳,+5��9dW
�E�P�EP�U�WĈ;D)��l,��nS�EX}��aJ�ZJ��Tc�����\K`�3>HD�@��E����Ɂ�^)D����x!Zm���q�𞝈r8 �����B�nP�Z����,�I"��� I���U��<���N!KqB���SY�������� @��6<���E�� ��^�����VxM@�G�jq��9�āW}�{���,Yf�Vd{4X]ь;"
T�\�(*E���?-�@�s~�,V�����,9mGAn&��(�UEIY�����Y�vfԒ4
�|��oƅ����eIb8H��¢	�p�0����`�ZqKEoiƴ(#�[�P��ϗ��e��A���.� dʲz�����፞�3�%G����r�gǬ��bh�yt8�R���F�V<�
�@���En���Hĳ0�����Ywb�b��GMn5p�RC��dd4�Y��$B��rq.|n�K�/�2�
�� �8Y5��"�lV��d��{�s�B�0x>�� C�,a��K���1����
�����E��IEH_Nzg���.����b7�5f|�?m�^��n�d��b����W��q�v�(�Ω���1�V(�^;Y;bccQ%�@�u�fW�T;�v~O!��*^�lD1���!�TJ�~�� ��摗uN9 �+
^)�-��B8�S��T�0�����8��6SU�;y芟5!�a؝.x��@S�QV��L�-"
�

Ir	؜�,E�\N�șR�^r���Q,֤�JJ%,Ui`�8���
fX=�.� VMi�Ç���w�m1h�aܰ����1���84QB�Chz�c��Ŵ���K�GBl|~�%�� wUv��7�_v`���3U� �a@��E�
��,4���)UY��[�%������%���w۟�S�F4��d�1��w/~>�°&!ʯ�)�y/��T�W$��!�;��l�����=����x#*D;p��l�{
�WLA��V<��N<vo\9*�������n'���m�j\)�D3�-�J�r�0fLu�C�euWM	q�D�B��Îe���t�M⾐s ���()B��_Ʌ�����`��u�~@v�p�F�8?���	����F��Jl��u_������ϻ�骓X�t�
7�M�iYb�?������a�kϠq2��$D�!��� �}�dWn���t���7�Ѩ�y����E;�y��EeK�"F����|&�N��'�2��0C��fY��B �P�����X�����jX��wtz�.8�砟���Q�6%(C�H�F�M��1"�ŅP����80��4|5�-N�00��5�v4�W�Zj+|�� ��}���Z�g������ı"	~���@$(��{�(^{�-Z��ؑ�����K$���3d�cd����6#����i��倡/<��7CF|��X4m�Þ�A�xb�WP�D���O�6h|+��W(�p�՗�⦚@�^�#�H��CŊNp�
�'�%�x�ջ�y/��;+� �ŏ����V��	�!W�A�D'>x;����a�����-&VI�S[%v��b�b6� �,�.aE>Kgc�,c��A�_��o��8���K8��,�O���CX>�N����1	I�����������l�j���д��7ǰৃ��*�X �6IE���x�#��>s/�+�jg���شu?gb�,x�n��q���
bB-���D�1��Ag|�u:f~���6�˝+����ps�
��A��1�B-L|�l�y��	��#F.D�\�A0�������hy0x�R��p�Y�:��l$�|���{�ɗ�h�AԬV	s�ނ�Na��D�D���[�)(�e�II�X�p�ˋ�T�I1�s�B��m��,LO1�m��Wy$���ހ�cּťf���.��d�h3�q�DMg�J��N3���B�=���"��Cg� Uv�A��q/݅� P�$8�X0a�/ظ�(��ZX+�Ч���vR�ɦ)�/4��y*w��O��~���20k�T����6��H�y�� � o���G>ޜ�5�5o��g�`��?�L;ܼNA�uQ�tޙ�֦y`�;�Ψ��(;_~�	�v�+>��g�ʨ�Q5	��\���Y	7��wc�̧���6��\����~�;mʅu�GdN!r
��*�����e��ja�;�Κ9�*�"�f{
��L�OC�|����g��w�|sؽW̕�%�f�hz3�o�f�"��Ҋ��:Q�H�Xr)�E�X>�$��S�!��u��T0aP#��t?��v5���3a�a`�K�UD�_�hs��5���H
��,�ۇD!���y<=�g�~9�.�ۛ��E���' �Ն3g2�v2�>�Ʒ7��N���Ե��ޕ+�G�
���M7e5���Mj.?mZ4Ľw�@�x�D�ikp #��tB�$�g��V��^��
�r����[��Q/^���I���������Q
�x���P<���STMoVә݁��~����D3;M	>���:� D]a=G��L�&����o�r���`~<K���-�|7Hc�L,�W�k�`�#
���A�M��qmp����o`�������8�)>\r�mގ�BZ�����������-G��*2����>�t�����0���r.�!���kÞ��{�v�>��V�t��We@�B�T�F]�D�֩�W���7�bO����+p}���5�����2�(X�~�"�Џ�n����S�u��Wf���=��7��}�3�Z�U��)D�X�%����M�xuc}�? ��o��>�qp:y���)�JYZ".�j�X�~0�μb�ӹ0Av<�6Xc�S<9�V��בD=��P8}ʨ{��z���c�r%��2��f{F��Q ��Ϻ�ؘ�O���a����1��� ��q[��i��?=�����dx�{�oEy��>�Wۍ��  �D�5zMrb,�'1���!��bb,`T��(��Q��J�}o�m�5�f����f1�lr���{��/?vYk��{�Sښp��Ǡ[W��ѯ��աP�H$��=PC���\`!�t�2�b̩G��6�+_��uM�z퉨��z�ch�I4�X��-z�ի���sg��e�������b��f�Y�q����n}7�ѬőN7�[}5�LNf���d���٘�����3zcƓ�1��9��H�����8�'&�p�;��"�}���w���,��s���و�yD��lT�
 Huv
A�qw$m��{(dp��mb�)�V+J���9l���g&�܁����RVo�ō��"]KS`����pbpCj�h0ۖ��~�ukC\pǟ���Ǟ�\}����u���"�t���ڽ�\8�	�>�U$�	���������c�1�� �M�vܾ��Y�_>�M���>�L��� ᷼��2�2��ѳ��Z�i�/�-¡������'~�W��k�
خ:����%���X�`Z�w�Ǳ���}/���]�Љ�s����Of����������|�5�/�L;�j�����`�7i���f�8D�)�k7��+�}�1*bs�Vj>%ĢP��#S��'	XKo��afM���ч�{�ɟ�_�^�#h߷��A���CJqF1�Je��(�Zгk0ᢃ�ry�_�0m����G�\����S��bA��w$v����N39�j��f7`�I����ѵ�Ud}`}+�����ݹ˰^�AU2�[���p�	?�N;*��������}
�]�~;����{	���mo����c�	;�Gf�/��G�����L�:��ޛ�O��v��S͆�p�ч��ú�*4n ���	��fu7�;ءg~}t?<��\|�,#�	a9/�	�.�궫�}#\A�`���B�sS�E[�& �H���JIP�m���`l�v߸M�z��^��-%
$j-�R~{#�����:#W���,�N99�M^s��$�V~��c�S�(����Ba�n9�B!��]%����L��B��j�Վ�ֶFxe6+� ��Ч_����-L�d��e8��ݽ+��V��oB}C'�c	��[��Z�e�䠐P��A�J�V�mCn�h�&���_��J����:\e��",听�C{فG�	�w,Q PmG��E���A��p��X"H��E#z�J ҜiT���d���ɷ�:��ߝ��wf���mM��H��ٔ�*�3E��@�z/�4�vL�ep#�74��H�P�\�^��"րnZ(�J�c����h!�%O����8�b	�W���V�%�h��ajUx�e�ښb���2m>���t3&���Dܹҏ���X�d;��x9�c&JtR��(����F�YJK�P�G:��lG��!���x�$�fR�|�ݲ���	��	����Qj�p����'��L-E�dmR�$U�n��1���1&�ҁ���>���9�����y�d��$-�N�+'acȴt��dWA�-�mn����
3���G6�!�Ƅ��#l(�uUӰ'ס�x��v�|*|�Y�ܶQ�J�S�6�@��]O�4x��\�\l���<�I�7��䁍�z�dP`K��""�<Kn<�<bF�ؒ���U:���(�]L��T*�#�E�"�� �]S^�	�� �u<(� 33e�Q*�?C�1Q�d[M�s���!�������7�CH~��e"��7آ	-����W�oƶI�-��!��u��x>�)�f����6TgMԷ�	9I�o���p=f� It���/�1��K�G�[3\yR��!�nh0��O~��9��Z䒭X,J��m0����.�E�%�տ����!,g�f��R�@��-@gG�qHt���'�uHPY'��Qd�P���E�;���|^f�cJj%�M��tb��N�,��QN�^�ȖCՂF�1�kW���c|��h�j�(R���K%��ǶL�t״b(]xAI���'���Ϫ��L�$�.�\oe1Z�IV@Wz�P��u�✘|�i(���h+�$C9�	![y��W��1C�AQX~Y�wT[�ZaHU�DL�e'��t����d�"D@6>Qi$�9���Ǫ7�D2[�Q"��V"�A�U2��䁂��#V����y
�<	�0p��3�U0c�eP	 ��ј�R!/*ER\:@�'˂K{�h+�u������|f&�|ɖk�)�>�_C/������!���	S�±SR"��v)'�1W�c�O&�-����8�����)�D&f_6�B�3����(���#H�g\1�q;�4e4��T !z\�.ȶ��ݾ��:L�$�/R�N�W*"��(�����tH\���ֶP��4D�e��W��u(�T��ĉ%%��R �%��c��]Au�A"��b�E�ku�ĥ
ZK�����\}+�C$j�F�at ;Y�t��/���FC�����nG�ן�~���Q�Z�+��. ��z b��5;���Ү*>�~A�V]?�=IU1�s\d�H�e���e�2���B�g�@	����6����L��;�z�=�tx������.���%[ذu9rm+�Y�����(R=?��J�Z���1��}7�2Pg�%C�l����X��2�f�`��T��mҷ%D�+�E���kuEu׾(���ld��I	�-�L��.A�V؊��M5��{������P0�P�g����ڜ9Њ�Q��,�
ꊆ(�_`�`����m��&��D��bB����R���>\h�*l��P�{ �e�%@Ls��rff��/�EˬH���ƀ(N�DgY�`x����]8=�����Ku�G�9W�e���p��b+��J����1P΋X�D��=����s�bS��?O���@1�������2�����S��/ zFv7`w�@c����z����8��?�4�1�W���G	�s�E�O!Ձ���$Y��I���f�E!�p��Opc���Q(�b�LԘEH%9J��1c|zǿ!cXAU�&|6����cp��=�d��|�vL1�\W���$V�g1v�8�<���?�F���ܷ�P��<�|�ƣ�g�8%�(f9єU|S8�=ޞw��{s�ԋ�q�Y�b]P���!08����8:mh�x���q�Ǡ�*�|�m%S���W��e#!�SO?�O�n�.GCeyƓp핑r$�"��,v����G�+�����{�$z=pᖋ0l���'^�����Q�E�Q��fɑ\��������gb�������
��I���S%-�G#k�����%M�v�c����T�� 4���cף)B�JIԇ-�=����5�*%��h-�u�E�`�Iا�g���b��y��ȼ�I���/�N��A��P�네3�����������1��?�� jw)�(k��m��%�$^�KL��"{��)�,��z��~�~V�}z9M8﷿��0bP��,�T�B�d&�1��'��7-���+����Z��.٤�N/�ӗ�Ð�&��ݱ�9��C�84NwI �4�\WP�0�x�Y��4���9��i>0��5u�$^Z>k^y��]/L�
�U�]���CA���j|2n�n*���.��H����2��C�ƽU��i�!l&#s��K�<ߚ���s}y5޻uι�D�kI��ܒ~ԨL813m�/�!�<�*�=a,�>��Df��������ܗ����0��?������JA554���o�|�<��d:������mH����t
۰���7��O��� �BG��XX��bP���G���K��㗗b}P'��m��˷�������0(���c����������%'�(=�׏���=�qH$�N��P4ѫ�����������a�%�����A��(��TU>�|>n��A�7�����#ű)]�(橮$��-iW?�cx��ؕlm`P���	W��O�A�v�
[�8�}��b��n��n�N=�bl�a���@ul��ٝ��r3
_��E3�Ľ���sr�^!�G�w��C�������ć^��LC#:��'�&�Ð�7�?V̺=�\z�)(�R�G�l��lT��-<��ۘ��~z�zW�%�a(PL��b�[�`P|.<�h��,J�{��x(�B�(�D�������c���E:H�d�����!j�,r�����'�����Y٥2�i$( k)�Y5�v��.ĵ�c�K�Z�f��y��F�
�CK2�nz��Ç.���}+F��U�o0{�8�̟���n�R��J0d�� _,�w#��N'�n�]���/���o=����.����U`�&&
ӌ�+���G�c�3��Yw�I�8�F2։K`�Κ�[�Əu�O9^�����nR�������k�t�p	��C��rXF������=�]��8�!Α��L�GG��G���'I\z����W%��Yh�(0�Y�	nM�An��X��$<0c<�0#T���^�v��̆i��}�?����h:�esVS��9ͷ�C7<t���;:[#���训�[�/A�6zVs���8��#��T�$�d\�m��9+����a��[�&8̒�@�'�d��g�c�돠W�ZQ���O����a���L�T��M�7�1�tkD��*�0c4|���h��%���E�n�-�uM����$%��A����v'��Xl(שVT�(߅��]w1���W����@)��g9P�!+.�Xt]l4�6]    IDATZ�G���=�d������	�*0���#��N��$!8w�]" 0��eőI�֬�2����"�r�g¢=�f��Q��#2�n�|�@���N�2��倷��ӈ8GC9"���'���7ջ��(������>���� �44��$c0�G�Mōl��z�����J�1����)��7�OF�{��K�
�*oL�����
)��j���������(��B�́[���/_�抗p����e�2��t�n�$�NSs
�W�ÂFk��߯G"�Q���-�d`�m������Nئ��BlM 5�RZ=p�$�����Y�A܇l� �=�Jl. %��g?W*r���#2Sƍ�2�ok�:�RcL��Y
������P�{u�D�^�\@��2u���y��w�ᱏW*;�$qL�����}/B�d5�$���u]��P�6,}{Z?z��6(�]`(�;Ճ7�1���h��Q�Ff���Z�c�;c'�K��!�٪(d���1[pc�����o���6�S.C[�V�y`�-�-x������
Ze�*�@^�� =��ɮ��kZp�3��ЩhM��zEށ�HW<X�>[S�B2��!c�K�A�o��Eӊ�� �E�/���t=n4�|�|5�C]�@mЪ2�_���xE�>c�I`�.�V/����tc`p���uT��X��T9JPhS�+Jn3d�o��p�a�?���Z�h�Dƽ���Z�a��b��|�8��\��v��.r#�IUk�������C�þ�C�슂�XJ,�J�+X��x��?�����f�!��F�k�1|�]x��T��pK�:�)_)V7k�.�:̾��ck����G�Qbjō�sN$%}tbYj/O�	�l��$1� �Wc���W��lW[T����Ӓ1����(ql��0m�?̞�k�#hһ�d�Na�Д��1mt�rX��$���� �m�K=u7A�T`��AWs�C���c$0Ȱ־؆%c�k:�H��'$AL.-�?�dZ��+K�/{<����U���E8p�uh��Q�و⁰]�`nn�_��������7�U3g
�W�0�V.o���ߏ�gޏb��pEԅŪjUU��L����%Ό��_�Y�������F��hYf��c_�b�fg���eH�t |���\�X��3��KX����%RXE��'��(�U���$�%�e��֎%o݃���_6Z�o)c��<J��NR'>Da�:������-6�O={)ӤӵHʜg�{�rM��xa�R<��2|�x�h�ȋ|�rT��@������Ϸ������\ps?�M�!V�FkW�1�ҩt�d�v 9z"��Y�$,����l�J:[C8����������|�΃�=�.<� 	���M�h���!�!����K��c+qȹ�Ь�6v[��6�翈�/܊�R���U���I��r ���&��L��
C�ƣZ�ہQ)>�gq��}��{�}\\��#z*0��c�o�c�D'���*��V�]���7���'W�a�eW�)c2ǨC�
��o�\�����G�dZk$$0�����}�Ԯp�}*cc`�(��O�1�&|8�5����'��Y`l�^!v��o��Q�Q}��c�;ӱK�s?y�L.��SGh%0���3�%0z���=�Dʄ�oC2F�(QNӢ�-���}����r~�!d�v���^�"5A��*��%�����*cl)0��І%o�������of=�]b���S��S��.���&Vn���-#�g�X���^�μ�F�ZLىs���$;�%,z�VL����ƈ�π�-�-����vu#.���{xc`���f<�X\	.�v�0|[`�;���E�?��x��r�hp���ܩ������Ģj�x�k<�\#�=��#�(Q`]���7����W�A�ƨ����/��ƚ��(r�ChO@��*���/+̐�f�(08����qS���?[|n���]"-�h�!����(����ͬ�%1眰?b�n�$ ���R���T��*O����ԂCϾ{��0�!���ƌq����I`DXN����5\|�r�	�"��� �U����c����jծ�WG��q�TsW���x�Q�nǏA͎Rn]�Ս6!d%����G��g����sc�*����yMܮFʽ�I4�����7�`���C���f��l\.�L8 �0w>�~9�A'AZ�vՐ�j�YƂ����g�boh��"x��U5�㢫H�.k�x���x��=�FlM��Kl�.]I-T`,~~n��<���;�!s	�j�F����hn*���f [����*��H��H�[�0�%wt0clu`���u˥���׮��
�D�@i���Φ
�@����	c�;��D��Q&G�z�Da���������̀p8�D���� �L����P���^8`��X��;aœ�������q�0�E����J5��X*:)�X(�}�tv��H�]a�`�� +�8u�,���ͺ(m��nQ�{8	"A��ϙ[9Qt=��8=!:�$o3؜@C����YX����(T f��m:x=��*��C�`uƐKF��[��U����&�Lc����P���1<�!���|�yԖV��)�����Ñ��Ќ�4�0D�����}�DJ1�`�̳Ǣ��Q��"<V�q��d>���.���OM��i7�*ge�,�]�����cq���LL������bu��0�sՈ�4b�<"�6`��5}�+Ǝ���%]�D%���2�MA4���<�����Ϯ�t�d�Ő/;���JҘ���(��Pn�n[���^@X���iZ�(�C�z'`�ð���G:��lR�}�cA�xi���c���&�8�%J|��.Ǽ�1X�eW$,�FW�>�N�]	Q�X_P,(����C����FW����/��'���iׇ�,S����1�D!���:�3�^��'\���{��ɹ,&wT�R�x+��WON���7���&Q�m|�Es������[31m�+8l��X�s���+�	��t�f��wr�?��7ހ�����7��6��$P٘��s�˜����[�5�����<�q�bէ/!\�
���2.��8
W[e��{ �F��W?���b�翇"���)nw	��׌`�{�������"�N����^�!���������и�<���06X=�JMXW�*2��i���d�E��[�]%����s-~w���>��0�O�N�-Sp��G^	?DU���`�IW��;�:���g���!��ފ���wb��7
�U��h2P	7��ƛo���z��=��t����Y6���d:�����B��R����:�nM�|Y��1L�Y��4��^��F�b�������ki4��+�_<�i׏j �°�
�Vf@9ЌLC�$�>�&^��{��9(�c�-M��@��_��z�VL��F$��rW"Z>r"I�$�S@��͝����C.{��9��_!��5�%�a�n(.���YcL��#r�[�J�x��
sf܌���$O'1���Җ��%��ō 邇sG^��']��n0�<i�-�Z�Q����]�}�nL�~���hW�5*�c���)+���x=��>���]ap�	��j��Q�7���h]��p�h$l�|^p����@��`Oa"``<�>X����^�f�q�\� �]#��x���9o�<�\{�Ŝ�tX1d�98���� �g������
{��TC�E�s%�"��E�1wL�Ն+�!&��`��D}J+-`���q��ǰ��I�$���hZ�0�Wծ�����gv�͗oY�sk�:�NF>��z��ȁ8���D�F7
��ȵ-�����$�<�Jl�eH���+��LS.\��
2(�x�w30�c��K��z��2�$*q�iZxc�'x�Y8�;�����?d��P����P���/x7����F�����`ծ�M�l���䳘��Z�s��h	����h��^��z��(~����r�6�P"�1���J98Ҷ�¾��ԛxc���q6�<e+!�L�N��O�[��>:�M�*��R�n�w����Z���/>����u�DdR��Xr�P�&�3c`H�U��]I4��Q�52��׺M��;��z�B�{��r�>��
�F�1�k��/F����(��7����OF;r+>��Oލߏ�f9#P>���� 
1z=��{}�'��9�;���e��� �8t��zvγhZ�.��L� �`(-�1p�LN�3�^���Vf1��ñ���G$��47���_�	w�L\s���͍�M��x2&�~>��GJ#q'	����xk~��rZ�*xvJ�	nbƬ
3pW���L���nAJ��&��h\��|���O>��w=�C/���ZvJ
Ve[�D�,,�EeC��H|�ٻƏ�ѹg������?P�ٚ� ��m�g�4/�P��\�7��*��h�����w�����"����5��kHy�W~��OL�,@9A�0�s�����
�ͦt�{�~9�5ZY���PS�;�e�9����y�)�
�z\�i*쳍>W��ό������3�E�������O��Âw_D~�Ӏ������Y#�+�wJ>k�w���Yhu�(�D��`��D�5_�GJ,>�AQ�d�.�]�l�M�����7!��A�>?$mG���䐋-�V���W�(��_�PfI1�*1']5"�Q �ݪ�!w�SP�����p�6X�Cw�$C+�JǮD�v��m��I&�Id�:x�S#=O�O��LCa���3(�����Př:��� $7��L:-w�'��������H��ڡ��dh&��� �K�X�{ ���q� cA�A��,�X��6Ӣ��+߈r�(礫���RS���&
�r��%��V�u������T8��3�>F�Av%�]ݚ�PMlK��s\�E�vQq��"G4?�c��Z93%�����dh�	�D:�t!��%�>DBHɂ��Z
�h,�(g����F�r�f4Zbmn�'{J\��4	�ȅ��
�h9+%�9&��X�j�S�G�\D�C�D�R�VY��5���j�*�[�(MPC�5��,^U1�4�*���G�Q��5=JF��O��K���HoDv����F����N�����KYT)Zn��ۡ��QZ���O��dq�)T�@���``�W�GR�\`ZaF�!'KD2�7�!��vI�óU<\I�*?4:-Ẁ%EYC��5��*Spefǉ!� �d
�� s��nW���Vv&JF��7C��L��>8�si���wM�2�4آ����
��+�X4VG&�Id�DEHyK��B_�B�b�A�N�&|<���qc�lή�a�8N��LJ�GE֖�O8J∁$fp*�q��񆋰�����	�;(F�h����E�1A?�5��Qe&U�(?CYw30x+6mJ���r+��H9Ϡ���d��qE��d@�x�"'�x�����H�Ӕh
	?�A�h�G?V>,q���SX�>W0��uTΚ�<�"j���=l�"J1�;"Pi��cgS`��K��e�q�O�9�w����羇r��^�p���E���+�n��7F��se,���QN�܍��<�B�r� ଟ�H\�g��cD�YX���� �y3U`��T�/t��&�b�RA+�e�j����<���Zo���yLX�|<.D[e�d�<�|���`�̈M�q�������J�F�|VTT�#Z���f��k,�~����U�%�kb���_��F�0�Y�D�v'�:Jd���?0$��jW���RW��M�'ʶ|���QGwm'���L))FUᤊS>J�J�C9�#�J��O�T]��U}Q+N��h��Ŧ��V���C*GG�1(���a�5��H��V��,<�� r��p�$yE�"_�~��<�f/Z�c_�1R	�cS��UQ-���QD}~n����/T楊�P��7�j5_��m�*>͍��%0�]��0o�|*K�
kL.Nt!7��Q�D\L�F��H-��,�<~ʏ����0��i���>E�x��,R�Qe����Ճ�o��0��]P*�D��v�v�8:�虁�T&=<�:\I&(}�YI%}Nf
�xx|H���[&��F+1:�YC*�Q�I�-�3k ��{��M���T���Mq7EƔ��*G�a�{D�I�ԋ�Ht�5�>�L��2~�k�i�fy���_���$z� Fda%$ y��gy�� WD@9R"־ �&�|�����B.x�RE���UlO�K��At�J9e>i��������.���{�*y�6�n\Ή�w���@��ZW܊����}��V�P}$�I^f&Փ�5��B6�Fbv$�������fS�j,�U sr��ḷ@�����"e�����ˢS�g�L�U�*���Z�!hפ���x�'���o"�m�#	��ƿ���N�W7����sjE�&�6�+ ��_Ԏ�8�����eJ��w!�	Ӷ�泈9Ԩ����F����rY%���!G��g.<7�H>�eU��p�u���:M��d�Q����S�CPwӎǐ)����e����ԓĖ��\����J�@��N"��Fw�جZc��0�(����%�^�Ϩے���Q�]�Q�ߩ ��3T'�^�����p��ZLJ�D�+����~��ˎ� Gn���:z	E������)�;��<0�4"����e�w��=�PB])�����/�p�У�gY	����ؘ+�q��P#E'���E*���2��)����Z?�[1�G�"�T��ȕJ(���;�QA���$� vٓ��O���,��*�b�Y������ి�WZ�ddN���rQ���ř��9Q��/X�Yp��y��ٕZf������k�����W
08�|)�):P<�|T�.�&l~��e,����}�y�:t�ɟw c�$�I���r��(zE��h��PcI��>)�Y ��E8�����l�[�s#6��b>+j8��EN�"pRhn/"��H�yT[�ީ�Y�n�RI�VR���� ��D�4��"h]���!i���e_d�S19��t�o%�C=z��rU�0Ljp� �����D|U�ln� �K�А��r������m�U��j������P����t+F�(q�e��P��ކOo?==����)�30�L�q�ЋT`�G��,ʬ���վeb������m�ߦ~����5��D��jt�H��֮Z�uO�n������) Ā ��/��^�\��;��mR3p�W���� ����ߧ�~���g����? ^���m	��~:����g'���=��hhk�@=�a���3b�Ӊ��bI����{�V�dQ(f�b�����؄��
�$ߑ?W6V;���S>����IU��to|�2 �!t�<ЬYX�q�������a�n�h�s�8��-�ŷ���wJ`���<�̟�}��?�;�E\s�0�n�I4���E�[����?c82f-��.C�����᧣*��!�=����m����Ћ�AZ�F,,�����нk�,�x\P��ؒ�0��I���@�'bz�O']�a瞈���F�Ǜ@�=��6�K�n�Cp�1Hl��}GIOS����X�(ss�|ci�r�Hؾ���~�Ѯ���Yx�F^ ��TZ�ʤwk����r:.��P󞲡8V&*�]TQ�4\ɦ�N}ae�0kҘ�)��w��n!0=r���7F,Z�t���q|�.~M�&c�u� ȳk�P`�Ӱ��9��F_�Ç_�l�;��E�;�q��Q*)�5�I���_���u9\5�&0�jd���i|t�Y���PW�I::'��J���>���$h�,���]�\w�Ht��M�b�]�_b��%�c�� �Ͼ�Z5���^JY�F��m����o<�`��$������b.�,�D��ǯ�АB3*Z��T��D���Qc\v-���<�Ja��F��^����)�H _n    IDAT��r`L��5���>A2�Fw*��qѡ4�,¦�X��͘���ÆǳMv:V�p��q8�?�9�-K���`�b2�v�w�"eؖ�ōy���Sq��k��o@����[~��:]z�Tn��}�]Ӏߎ��G��t��Pk���� C@��q���SC� di�(]�����.����D�Aڬ���E~ ��5���%T�!�~�6r+���N{��������R�t)�#E���������V�r!Tn��a5_2�ć@=M�\u�����-���F����愑�S�{�g�����.�7md��Hī��K��c���q����2� N��� vqc��D2�hKl��_�p��I��9���N,��0e�p�Tr�MXo�@�܌�������.]�t3��Db�,�4g��=~<���V����N�M�G�.�jmz�5�� ��8{�x:�7(��mV'��!�r¶��J
��KRp�9|3�֭��CQ"�?g7#�P����;	�������h��uߴ�Wˍ��7����۰��u(��%> l�"��D��a��/��g��]�O?f���>i�w%��y���G]��!�!��'5�$P�*���UBn�L�|�6<x��02=A���t��l��އ�-�Ѽ�+�߹��*O)�8+U�|����a�~�$6��	��[���ᦫ���[7�+(�H��bX1\x���w��ж��b��y6n�r(���	ߧ1�����A1���+nĮ�ׯ���j�2�L8�kg"�5U(b�ϡв;>.�n���Y�W��+���X<���+�Ҏ�,�Xl��L��r���"�Y�f��?F�b�YW2l����n���-v%*0���!N�zԉ���q]"A��0���oc��ɸ��+��-]�h�h)��e�q��p���b�����c�_oÌG���#�K%MGm"�EkҸ��;p�W�X�z~>��t�t݅���C2'��o���bI�2l�����:��bָ���G��s��� ��I�z�F\�}~zܮ��uF.�e6!$��إ5�c��O!�Ҍ��OKD��h�(��j�*���\���d
���o���h��� Q�r����2w&�\�O+�O�Ƞ}��h��)�I��w�<�}��1z���.>�}��]��z�A$��q�H�W��Ϟ�.*2J���N�c<�i�c�U7��F���B�j)>Ǐ��,Kj�`�r	�(����f�q�yi�q����O#ѩKW��p���i� �sɕr��ﳏ�-�<�R�r�p��7.#���������O|�Q0z�\�rNg���'��U�6�a��#�܂���	\����Z�݋�W�[�"��ʪ��q+�cK��nį�*"�c�U�SE��V8�72Ȭ���9�c��k7|�?���I���rƘ��މFԋ�,�Ǧ�"�r�x��JM�.��#��[P�P,p���C[��ܯ��?%��r�V|��A�vqF��[HB|��$v�y$7�(|��k�uie���+kh��;}���;�K������y��CUu��Q�.�:C<��y�=���Z]_R�������wV��'̰��ȥS]����E�����%�F��j,�\"��R�������޶�����T�&E�BU�wZ��d`�H��ȭ~k�|�A�ƉM��m��Ʊ�w�	�;�1�~75r:�|������ yq�!��2c�+^X��S� ��a`O��� ����^�h@f���*rT�*�����������Wym��y�op����g��9�Y��O��M:��[�Z���E�^��lK�r
z�,��U�R䏋�����Q��i��ŕt���
�韼8W�Qo@$u����|���H�iV����nD���ĳ�&�u���{�{��3G���>L�F���y|���(~�*Pj�11��!��Ӱi_�`#��T���-�~$��L8�ݨ�Z�ԱPR���M�'��'�X��^v���d_��~������y2�R�sz��w<���*4y5HF�'ї�3c00x����g(j��J`Tgj$��Ѱٗo�P��e��E����^S�6z�S0����QQ��MT�mȯ~Ec�97#n���1��1e�#�9���O��A��ڰ+ߞ�?[U,Tn�T=j��p��1Me�
Eo�����4��=A��Wc��z�	eSs$�V,�D�5V󏲌���B�ΫG�lu�������5?G�
:g��n:��Gl
��<���D_G}؎��@������V�By?ɵvEZR�6��Q[l�eC�yM�Q;r�ȕ�����A2�����&�FJ�^Ɗ/?��a��1C̾�ܶ;o}����E�����!QX���ߏ5��EP���iM��$�@��ʲ�B*7K	H�/b�*�XL���h���h-�D�1sk+.F�d�O�	������E�1�����U�4A����@��� �_�ɒ��A�09J*�d����5��ϐ�E5�ڕT��Y9"3G*Ҳ��M7D��:rR�����_�
C��b�QGö��$r<ʨF��D�I7=���hcq��j��ȶ���ӑ�[P\�*V~�)vv�pwgO�6��Qm�]�z�?;����s�9J�%袷c��w������J�<*�Y�������Xe���:z��#�n��Q2Q��+�o}��n�6
�Ejn������=O�f��@����y�}������������<
%t��a�p���"7�j|^q�L	��M�TA��(�@(��O�Q,{����d09�Y�T�������!(;ΐ+�2}1���.j�k�Q*����]Wl?.�X+;J�Q�GU��.i�"��-���s�~�8�u�(�)�F��vu�O�쬋�v�᷋!
U��X��d4}� _Ā~c���&����6\Q`D ���S�CJUc�������lt�AfxCd���lW��d�=���D w�C��r�(�[ø@�C%�O{��Eo܄���hZ�ɺ8R5�ZĬ�̅ׯ@�ϡK���)heq-@�m��M�Wա�~�~��W."nSۣ���Ĝ�VJ���!�������wb�"a�!��]	��î��������#�=�-0: ZDj&���.��$� LG��Am*���q�b�N]�u�V!$.��G6ׂ�_D�>}Pv������epةK7؉*�3��H!�H+�ǆ�b'KvB5�g��e̱���H`�}�Ň�s�o���Q��|[`t<c���bNc�%e�+-&Qd6t��$@�Z��������%�;%�HQ�\C�i���	͙ft���U-{�L����X5R��a�q�n ǈڬض��ص=`�ꐰ���,il��2ƶ����EdbQ�J,#0���D��Cw������"��:��>GU�ӱ�f�R�.Q�9��T�����k_J<��g�y�X��ֵrĕ2^�K<U��E�L9'lE`�O�e�!g�~ʗ�2��Vc��͔9��3�	����ۑ͵�h�[�ż7���K�h\���z����~{b�;!,瑬������,�[odJ@]�t0�^��b��ڶe�'�5�K�2�$ I[� � ]�t���X`L���qC/���m5FGj��<�E�̒#@!�Ќ\a�����n@��yX7�E��i��ð��H8:���!t��HR RH��X�f-&M��Oޞ�Ԡ�ѵ��j5XղN�
U��H�k�20ȋX����-0Tq�q��NWB7���(#�s��mhA3��%�
��ڴޒ/D���}1��Y��t�2��k�����r��q7�/~Hv�vA��.Ы�Qݝ;���Ȓs
>�f%�q����e�m�gǋO.����Lő˷�n��Bz����n��/�Ev���i���'�
z�ҥO?���Ԇ6<�G2a�-�ʮ��;'ބ��yI��v�%�k֖�������+Jb�ǀ�ʐ�FB��hJH��]|n��{��� ���|#�$��!��)�cݢYh�`�;dw|��,����pvۡ�?�ڮp�	����T�
�n��?�$vؾR�:|>ov�7�7����a��G�h�@10�1������Q񹱘�B`�5~���uҜm���T|���	
�X�~B��TM
u5lw=�~�~@[#׎�{�C*Y��m/u,Y�5vݥ?�|��;�X,�;n��=�,RH�-��yTW�b��ň�vG[����T�G��i}�X-��pI�)nޕ(��p�o��]��G�F��j�ge^�Ѻ�t�3�塃1�曰]����j`��siT�m̝?��&M��rp�mwcƣO���3�V�/+ee��_�#~zjz����?�����������I`P��(|%I��%0��ķ��ಋ�������V��^�����57��Q��in��ӧ��v���HC�|�,�f.~pȁ�a���6�A���V<7���\Ĭ �����W�m(���OD��' ^������D���@qy�T���1��Vo��X�+=�G"��^3kg?���<�r	5	wO������N�z������KX��B���ؿ� �KG�/�tt,\����wO��{�~�����p��GB�h"@Ae��E������Ə>d�5ƶ��x`��:a��Cqo=V}�:���b��W��n��X2Ҿs��x��ѣWOh�rՏ��4��B/�Ìk�X�p!v8wO�S���୆�_zS&>��G�����^#��[�%���m��q����U2��p�lW��liٴ]�pj�N�
��2Bz�S���Q��aeW`��᷿����XP��a� ��q�ģ�>���	a����!�l���F�f�B��q�u�4�$R(�6(�����e0�������Ъu������U'W�1�*�@b;h ��G����[F�ő�^�Px���j-��x��G"��.>�z^��L[+�f�&���r��FM����^���g��]+�懯�	R��*�m���ǟG���#��R��8�X�r%z����M'\����Q*�D�xyc�=�|�8�8��;�A,=�T���j�AJ�	P�N����0=jpu,0�L{�ء����H��fx��<�Za/DÇW.��ϡ�����FQhCJˢ�q��S��:)GC>O��j�	�x��'0a���ڥ'�H ���͵��@{.��+W��_��]�r��N�8�l3庐�}�I{8���Q��1�[���U�db�*h�B�3�-*G�1�߄��,����,0HhA�=~��Q����S��tX����CY��y�V$�~�N8nW;�(���P%aHc���3q��Qߩ�D|�t�@L)_D"V/��_-���O�F�w�L;H.��6Z�"�l����n�8�0�Bہ%��}�H��|Z��f0����m��OP���y-?��~��D�n��$v�bl���X>���]�{o���&��ke��ʛ���?^�xʑ����#�+#��(��T��r��`���8�����s��%?@��{�K�>�8����5B�jS���QW���1���a�؏'�߱��=�=v̙#�=��(Q��{�Rr�)W�����ĳ*$�:(�tۑ^�!�~����}��-$�$f�������Zt�^��rG�������跣�a�FOk�҅M8o�i8��(��$F\5�8�~����6<�23���ZEE``���u�l�`>�;c�8�h�P�\�IA`�!R�
}]
t8�!SJ����k��_��d�r9�{W|��,\~����E}������NҶc�U��k���w�{��B���I�
� �+�b����8���p��g`]&��:����{�r,�2�vĲd,`�HuY�%��m��]��� ��A�;Օ�S`N�V\��22�Pη�q]��6-��~�4���#q���ѥ�u��#T%Y5�<�����ѩ7.9
󾚋;@�/H+L%�l:�5+��1c��1�'~]�9�H%��RH:5���h�
泂���w	�=*>�e��g�
J��t%�(a`�e��u6�'i�C�
i���
��кA)��d'����2������Q@���I��!��a��F�iL{�>���&��=࢑���/�`��v�C�PSǒ���u�n?<Zjg�M�����������V�0�-��7^|���S�}��]��N��9}�Y�2���n��V�;�'X�Q*`��X��X�L$�<J�s���;�`=�î���Ʀh-��࣏��Gg�b1�Z2�IT�m��W'au�Zlק�N6��Wd��G�.G��.��d�D	1xAA)�TT���d&"
;¹�-0��v�bJFd��� ќ��G`�f�+ۈ;&� �}V�{������4����+��@�����|Q�3J���I����,D�.�L{�k�d/��o�E�a��M��(+oڍ\0����C�S.����Y�F��\!)�%EAS�#�+m�����(���ˮ�QhDz�B俞+,> �g܃~�C!�G�U�l[;�S4��3����1삑X�p`uj��ǀ��%�h�+��U���f�N�� �[�wQ�����dE8j�P���Z�m!0�T,v�k_�Ppې).B�!Z�Y[�̪�X�����y眂�T́S�P.`;:��툧��vsXٴ�~_�nB�� x8�2y��6���n��B���6�]��١��������1Ó��2n��u*�l�9�SB*GG�U|n�+��E�L�$	�U�as�ihI�E[q9KC�n;A+���䱦1�� \C^�0{����llhX�҂�\y�qe���>���]Q�Q�Kؐ��"i��.]�"�̒XT(�f����&��VsW+�Q�v<0�+��+��E[��h:ׂl�
;�e��)Z�#,� �~|/-���6�X�0ӪtA�����F�^�D����Э��ր����iȕ��PLCגH�I��d��|^��
G��#c���Z����
�o���f�^�����@;j{ht.2�۾ȱ�c¥�L�J��mH��D��Z��8VI<泅"z��߷�[6
���7ÉU!����T���D6���DcLi&�"_-v'�B`�9�#RKӨ|�K���۽=b�+�v�7�9���T���*�"U���
�S��x"���FÅM�����~j��6�AP2���O�B�?yM�v?�Z�Aw �MP���3��110Zڰ�?�*�Q)�"��)4/5�Q)�b#�klx����;���v�hȣ{��0�N(�<z���s}t��Kp§VƲ��E��o��Q(�g�$Cp�B������9�)�U_���}�U��\}��8tQ)bP{ID��D����E# �t�b/4iV�I�����X��Ac56l�H?e�U_�����A�9ƛ���Խ�����o�D*4�����pp��;>[�s���ɬd��=�|��aL������Z'�F
��gغ�Q|��@�$p��t@�Z������lJ{�$�o�`P�l��P�l��'�B/:&��2-2��kCiᣳD[AFGb��o9`E��=����M]T��),��;u���g_���>�=EjbP���o��j-�w��0�[r�9�L�Q],#J��-����!����4GQ ���b	��B�RSW+�B8g�l�Z��ܹ3L3%FB�%~��i�02)�LR(%�wa۴ќ/���R2��:\TY6�n1��(}��%���kW�8�8���o�Ըtᴣ�H2���>y��e؈��2�I���O���~�[Q�4O��	q�h�)�+ތ�C�,������$�P�QsT�D$�P\\�pMPuȐV���S�9�����C5/�s�-�'R9��I��0ۨ553v3bR뛰z�cF,�{��vJ�7�XDb%������5���u"�I3T�E-ơ�_q�B٘���Js�ZE����AnڼA���:����P��#�!)�lK�hD
���ɩ�}!Zr    IDATj"��ޅak(� ���ס�<�v����F�c/!����7p��kP�ұr�؆�g�G�ye�<|�2��4B=�<������'� ��,4r���ي�Fi�JH��b��%>Q�{�LD��\C{��Nhs��n��NQ��X�r�[��1�\V�%���ka�E�b�'�iH�%��d9�>Ǎ^�sRB.���dV�#4��x�韢����	��nC�bT����Cc;�,�:c2�XS+!0QR��c���Ii�567H~��f�/"b���J�4j�E}�!2T����F�q��Q	A�sX�z��'��ٹ�lh��Z��nM?�yZ�?�������n���x����\0���#.|��y�`�d~��76i�1<T?ŧ�����X��3�C�V\,�Z�J�J֜�[�3W`Ř{� H�UIO*��Q�$HH��,A�����4ũe���:�*�'�YʑV���,v�s���p�5ȥ�F�q�/�7��I�T�7�ݧI�ք�π���0���Ȕ�"� �7�2!������	�u�X�3YqJl��V����6��L���s���Qc��7�q�K�2�48�V�4n��:���S�d�l}g4�}	��~�.�]:����?jX>��^z����{9�ҩ~;x�
1.�v�6c��?��g)Z�L�l;����u"���w����X��I�.Z,L�b�Bj�^��d&I�`�F�4a����Z����\1���Dah�G����D�����%�6�>�c��3М��J��[�y��4s�&��_�Za�%D��8��r�bK��bPI�Ee�C]���X�'?�&�y?�kN8@���0	��g��(|�7����'����"�����~=�{`%:����7�v�[8�2
5c�	�o��g�P<��M�بu����h�[x���h��v���J?���PY�#q	��Ɯ�%E�J�j�>:�.�.c/@"!�R��"��1�o�y�B�R��\/'�=���>�y���͘N�3����<�*lF���N���n�ZcU�2�A߃�*��GEf�al�S��]�*�`1A�B�)wV��$���/f࣠�R<j�J�ÒԆ�S��N���b��	�ϛ��	Җ
U|[�m��`������q��}kW����@mFów�m�a,}������Ѝ2RQ��#���PD�[? 6��C���,d�<����%��5��kV�԰��.�?��E�+�NW�X,�6-4=|��&T�7�ȁN��G�c�^]PW�UR��:	]�g�a�+o �Wo�U]�IYBF������Z%�#�Ym����kk��� ��л�~'��f���	�p8 υ�j���EMW��|T�5_��";�:�ݫ�nb���@�$��*���B���$��T�(8� �9���C�ք�����3�ǡ�:I��n��,�nC���}�p��*�}�uq�lT�����x֞=Ʋ?�FOX���/_&��je�Z	�pa��3"�׿�w���͞�Դ$l%��i��E�dS#���f���S���5����a�U��0(�+�S�j�ç[��>uN�t5�tG�yr�T,Zp�w��iQZ�q]rz�6�N���}6����񻅓1�4�ثtS����*\�pp�sp�)g��r��.؊p���a�O��6��w��
[����S�#�D�DAY����P-V|�(?��
 ��nI>U(�5p�����bOĤ&,�P�0$f4�]e�%+_�߆N�Vl�`%��9�׌������6WF*��>��^_�A��$�}�s\������|��vH>������4��G_~���
^	Y;�XD3D�����_nŃ�_�BQ1�f,�b���m.��q3N�trF-�������Λ-(���g����?ؐ���ޅ�_~���T���E�1o�$t�I#�Pq�D�lW����&_�#�}>r]C�����K0�dt�Tˡ��&�ob��M���N85}��Mn�Q%��|"�闔G0,9���(�K|���1ĵK�h�Q0e���p���H�n�H�͗C�*dZBHk�XT�_W�=t�Aa�:h��H�p��Ǣs]=r�2�ٯP�:�G��g�J|��5�q2v��n۰t�{6��~��.7�_w�FI�D�M3��<�a�5���g���y�����Y[��r�J�̽�;�Z4uȯ���~�hDl�H#)%Ib���ֺm��{pԴ�تף�^ċ7]��7�E����x�#]�@Oa��Y�u�w��_J�X}�E�oҵ[g��s���=�U�Kf-�~������{Ҍ��+��bpfE&q�
���5O��-[��E�D'����+Sb�J�a�e��l]���b|�{�y�'2Vb���f��H ��BQ�yL����	6��'�|ad`�����ա���oF������8h�I�_����ƍ�8��Eبգ�
�vP�-�P�|��>�w�0�Q+ՉC�t���j����믽�\v��m��-�_�1n�5J�V6l�#�"����<���n3mևu�E3^�w���.���$&�R�t���ԫ�����A���Î�xc�EXx�t��M�C]��G"�9��%8�ĳ��<
[�l�c��Z�J}��N�#<�[֭E�#� ��3��Vj��<��	�+��V��Vd�w�w�{�%C���B�t��;�e=�7�c6M�m�nwjPpT�>y���M^$t�/�~y��ym�J����GO���._��Z�f&Fa�=�ϡ�����"}�X�a�)��]T(��[p���PHw�֏V#������	pY:<^)�k60c�8|�4��BU،Wg_��s�a�n�%���d?�UDhW�҉W���磴�I�Z^�sn�=�;�*��I��N-.�6O=ѾG�!L�$�I�Q
)��X� nhH.�a�Q�t-:�_���q��:��FIr�\�l���Y�ɍ�E!��0!���L�72r�U\�-�e�����'� �����+(~�	����v���>��1q�Ͽ>n	���a����&�{mڀ��e|��p��W��K��b��YC�N�'N���hX�.�=s��8yW��-#�P�t�R;e.6k�P�f�2�GX|�4�����R�F=8n��3.�<�>���Kxe�0,�?��v�N�&�އ ]���N<��ǠĘ��(Q3�J�LA�(Sn�LW�����~��ʭ��3ɮ4R�@�XϬu\�C��r��%��]�N��Ft��sa���"%)*�3�JDۃ�?;�,�>��g�dt����m��.nC����'~8z��=�ipI�5�Z*4�4���M|�?����Q*�15���i���<��'8a�Ll�jѼ�cl�ۃ�9f(���S����G���|ڈ{ߏc'^�u��m��6�_�����W���^���0�;������(d5/�5WL��{�iS�̇�a�Rȕ"\y�:��{�-A5"�J4\y���K�xv˚�Z��m�6��P��˔�Th,,ɧ.#�$)��)ZN2"߳��+��
nYVa:*��4��_�(xe2��]jhȗ����ݭ����t|�<�]<v�e��l��۱a����c�;o�h5v'5A�YB�¯���3u�ƈ�(T�5o����/l>`nLшJ��{�V5fp������BԼ	o, h�8���
�2`UZ=z����m�[�_��f.����ZD����W�=c:|�l�PҪ����3t�غ8�Bd�
Bt*7��\4Y�$�F`š$�J4�����.��G� jvg�3�f�r'K��L��<�"�4;+�)n��?�5<RY[��v7����5,]0��=NW���������Ġ	J�^&8�q(��P���?����,� �˴�NJ $,�z
�Z�����Z^�]#5|F/������k��B��b��.e���]�^N~����2uxF
MZ�T-�ЭC嵫�5}��r�8t����G&�$qR03u��Z(�5p� �\�ݨ��ƘGY	X�|BW��=�X�rv(�L&����Z��bq���L
㲶����cIӦăI����a,�n���Jsg5��R�� mZ������%N�a���m�7������?z֥��=>x�]j�J�P)V+ ��z�$��5$Q�y�� ����N6ZaR����
�/!��?�S�%�)Z��$�/�B��n�(�l=]*
��tRI]G�L�͗$�Ϧ�'w{��1E,C,Sig�Q�Z>|*7�z��H�$ϰ�h�[BZg>	P�N�B��������\�<ߚ�;�bi�x��}$������?��vJ������l�ǃ5zv�2��)�ѫ��)��B�h3�q[�1��ѳFL�����!1�x���u�,Q�T:��H���2�ZYk0����"�mnCJ�0*+v|��\��i��Ȯg I$���d��'�?G�ȫ�	��l�0�x
(D�{.��O�0� 6o���J>�˼Df3>0���h���|�L����K��tV�	D4��PG�v�4ĄuM[��wx�7�F	�
��l�K>���x��sQSi6�dh�Y脍b+�_1dԨ����;�Y�c�d�Q�[�j��6����6�%�i2I���>X���y�]J[�P���q:L�Z����BX)n)�n�˓��SKOk���؅GZ-�/c|�|/�&O�f������\ض	�+��<���m�ek�^��h������j���吧�x�>ue��}ʿ4]YT	�21�c���'^��_٭a�}�#g��<���x�3���5�a��C0c�.��.<�n����)W@d�ҭ�}urwuch�,�q�Γ��U�R�N����=Rv_=q�K�X�R�`,'�a��
����t�e��'�g�Zm|@��fg	� =m��c4���z7�C�b��7%���6e��R0p�$��SQX�+r�R˴�|^�x��7_q☑C_ޭa����3FM���6F���-jq����<{VTF�U���&|�H*a~�'�8�e,�[&�q,��-����8F�!-��	W�Q#���"��ƀ��7QCU��)i�/�I�
x�~�s:�*oD�zH���?�c�����<��3�ﬅNT�����P��7[�<hV�
Me�����Z\��E�b����|6/[8�ї���=�#?5e�/�j�"�a�mM��r�FP�4�ӷ�C�k@�cI^ �c�ſ��������?���RS��h�x$�Lx�\ghе3IV�Q�;D�h1&bw`�=�1M=8���֎���o�m��""����@I�3'#��.�� ���vu�c1<��lGr�b� ��ѱ��p�K���!{3�2�7�+	��BI�1b��-[8��=�RQ������d_�Ca�f?����x��@����m�k�3�J�.����s *��{��VW���{�L�N	������x_>V��P֫��G��ʆeo����R񝯖������\8Z�oy����,r0�&�RA�mNUʛ	��cP��=����8�(J%��f5M1�7W���Ο{��R	1�1�'Ti�&��r8b��Cy�����,���*!P�,F�W@my^�c-�=��0�+��R�mj،��M�&O^e���a5�C��5S�'�T�?�\d�U(�K0���،�/���D)�/�����|�7^!�iIN�XLOb���n X{�� �I �A/lDgm+�����=������ҵ��0�/b�[����,�vVD�c����������{$��'ޗ�O�>Co��ϡ0m��C'�u�-�j���0���%m���w[C؆#WV��8�d�E�]dc՝�p���ثc��^� L�����T�|�t���2�F��'(c�c�<b��8z�5�g����!й�A�+&�1��b	l��3)W�򐽗�߈��F<s�L���Km���`��X����`R,�*���롇��F���;>r:�:�ރ�/�OY���%�jh1��;X�%��b���F������=��Q��������0BW��$�e�ni�q�=w"�u�W#h�{7P\>b�T4��Wk�P�� �7�6u���:�z!o�IBC҈S��\5��H|�Y�Ӵ�����0d�	�]���ų0n��8f`/^I��P�X8w>V����D�����a�3X�a�~ElT�qg�!L�@�h^�}\~��i'��0*�mhp�f[ҍ�i���7���5����a��I�֩C�W�E%��KF�P�9�N�����u���p264E�b��8b̵�W퍂Q�*$��\��R�������q��&���M!�`v�C�h3�_2cƟ�c�F�g#O���ebѼ�X��[r�bt����܇|DF�N 5���GLG�����`i���=��%܄�w��0dEqʜ'��1�&�0D��E���T�(,�3];w��^K��p���O��N���=dȉ�B	�����3�.�c���Y�����z�l�1�I�]�<ŗ5A���v�n����DegK(�d7�&�ml����7b�*���T��[��v��y�Gv%����2��l��X��s���1i���dInO���<�J����U���ѹs�j���	�K1BF{^C�R�95e��,��]�|�^(Y�`�Q��	A`�K*1-���~��8W%���zzVP����%31n�98f`_�0�"<±M,�{V�Z�89��'�{�=��c؈��}����,�P2
s���u�s(I<F�c�}}k���h�a��C	�1�4��蓙kT>���Fa�܉�Թ{�����/�a�㹫��x���t��]�u��rfM^��hJ��	�gF�d��c:"����� {Z��C�a�2�����lØ0�,;��pl�*��[�Pr�\�JA[ƞ��#>$a���
�_(�q=�8�������+���y���2rҼ?��0T��鞮sa9�,K)"������F`��ɨ��M<���ɰ)�#GUB	�4�{����O��KGHKPTL>s�O^�c/��l/�*��M�����KbY	��'&�_�0,;�\-;(���9�_<��� ��%M)��0eo���j�W�{��|.��JP��a#����ֆa��v{�6Ɗ�;y���j�a�a�^=�1T��:�1�\��2̝;]:u�K�{��#b�h�+WUɨxs��Æf�'-��/��L/A��&��$S@B$�e�QC��;��v�-ư��w� H�)2�j�~�B��w��/����$��m,�V�z'|U�=��r5f
����/��.إa�Y��QUI�p3V�qyn���C�8D��G�9b�ܧ�b��P���Y$WFd6�mF��1��l:�q:�Lnd���0��F��tT<���Y'�de�7��s�i8��d�@� �|��}L��z�8��ӽШU#G!�te�k�#LH�T�S�J8�a�T6���vu}��q'�9���L&��،��zl�3fa��q��_���EQ9�O�馛��悔ޝR(����~�1�8�7l�5t�$t?�:�z&FW*��8�!��k���RU$��p�%��vø���O9yޟ�j:�N@.��%�!�/n��gxeŵ����9EN�"L8p�Uh�7�?<�1Zݡ�^E�E�
A�AK�n��à��(,���	��&V��o8�G���(�(h\Z,�{5z�$�P���k��P�ʎ��ŋ)#QH+5ZQ�$��8�r#:�#8�6�����e@o�ۧ^PhZ��]�^�����o���JV~�μ&O�����=G �+W(��?��ngM��� ��p]�7$���{�kk�1�m���؉�L�����$� �M�8V��	�x��o��A�l����2'�B(�Co}:c�
�o�M��\����gJ��􀓿-]��⺃	�
ƺj�1QT����I�P#���![�c���H`}
�����l՛aI �Qqh�z�    IDAT���_��@�d�-\�����m~�GT���.D�Yu�Bz[��T[ �:�u��0k���|$�&���0�$�4/_4��=��v���q@�d�+`��}#ȣC*@��`��HBƜ���t��bHJevo�sۊM���Bj��mo���Dx�03Uȗ�l��I�0��I�������A'���+��Z��L�� /@п��U�CgF���/�1#�V�^!}�+P��x�3�*q�2�
~��c�^��A��Q$a��g	L��6�hv&n��}XE+�Ð�Wo"M�,�f���<�F"x��͟�,�ui�E)��ga!�D���#��,7�\��!�/�LjP�CGI))<]�O!?�0��&1 ������)gU���9�{镴r+���*A�:4M�\�҈i�g�[H�j�c|��j�ؾ��g�,����6?=!#W��Ie�FI<I��\i�q�;k�|��}��F�rAC�)� Nt�Q#Ur,ͤ��y��l��(��%7���![�fkP���?K�6�} �t�pG���2'�݌�܎������??	I�)����"�|aK�Q��G�c;!�8A�DȈ6;�b�x���R�>����+8"��{��q+v����x�$4
�z�X��uJm�6@������0ڄ�jWUR1{Ob�Z�Qw��{&�+�2d�c��I���Q.Tx���(V�� ?R	�Z�yTF�����.�X�����_p����l|4��7�#Ij�O;i�I�T1�ib�\�?5*{�X��%����0	K���(r΂iā��(�[b;3�؃%�n4.A��Z��\v�lE�m0�ۨ0���+�xbl�c(�yk��&�h_�+nq��i��#n)#����f�Ҫ%��!��̡x�=�:�L�S����Gy �V�^*���X̋k%��l�k�ZO��c=*wGMg����Crbe�!�8�I�+�Y�0i�'����sɼDȢ��Ğ�>1lz	~�xO��U��k�O�?!k���%��Da ^)`4y��z��%$w��hLP�x����7Oo�-q��J�t�+Hnl�	�I����O�ѿH-�<�J�8�����[��s���-�S~�1���l9^Ib���mx���-�ɱXFȄQ���v9ȚG쩨%ƽ?R�
���q�{'�xw�bj�4}al��"U����h|��]�֯����cH����ю骂ޫ�͆��bɆ$�'#n�8����$i����\kI�*�H������_�Ժ�3$V�5�0�¸�&�^�k8DV��	h4�c�v%�xr���Q8��p�̟a�+y�R��^J����7Y�ja:n�����!���M����r��GM�G|�$�k���oF{��u�j��Ee�-E� �zc���B0�`�Eۑ}ng�۟���M$y�� �a�?B���a�aҕ���G��� �Cl��&qd퉇��J��1q��i��ai�����~\�R�Dr8Z_�T9�G%{}�o��j �S���{�>Lؾ%�r��x�v ��tQ����j�I=%� C69 |H���sw������#_�8f2]�ױBH�[�Z�&�=.��	��!���7��"Yud���?�*�/���]hh�5�RQ8�T*\1�������D�5)��sԿT�Ί-��Q��ѹ�����i���%� Kj�4��%=^DR��� �Klb:�|���x�<I�J�h�{��H�2C��[��S1h��e�P��k@]M��7�(l�WjĖmM��J�lMg�k:	�g!�����0"�?[]]YH�]=$Uٴb⑊C}�@�Z!�X�������
ٶ}v����[�ў����D�/u3x
�z��E���!���FO�|�r��b-yF[�dL/�=���Q���lpe�r��|Ԛ6�}�W>|���V:=�b���PW��|�lY��"��s �p:����EIKAKנ�(p�>�5�@k�QM҇V}�=>�V_�ŃQ����`_��a���}G���2��˜C@0��|+�B�$S��M0��	>���J�RNO뤬-��g�B�LF#iH��뜩�ѻS5>~�oX� o�N�C�9��?2�(����T��o���<�L�|*`T��w�G�����ed����2wQ��˅�(UM���V���*��dUA	ͨ܄��%�b�P@�<�����ٴ��5�$g��)�+w�U����ln�)UwT>/G��IC�|�q���m�z
��ADb��ql�?��*-,�n8�����r�=��A/�?������Ko��OEV��hI`��#n�y�o��\���y	g�v.��0q��[���g`ejĚ*�q�h��jy�Ʉ6A�WtYHRO]��=(
�?�+Ir��*+I�e�̕�Lg�/���wa)�9�P�V���/.��'P���z�s�L�, �ƢIĮ���� r|R�U���^�f�\�V�JbFd�7�ؖN0INI*�5�%��n	�TVi#��>���/�A�{��A�^��|�����8J*���x�u��w�Mx��_��3�g�ES�F٠�ԅz�Xצ��LZh��*7��L̻U���DtԷ�[��͊m�u� s��?�.S�(f ������Yp�(e�~��$6%gUj��G�l��앴u���7Q��B�D����	�1�����q�_�~{w�
#Ij �8VUa�B|�������Kg!_u0rf�����_�� w�L�M9!ZT�_:��D���t�6���3p�����?�S@A�n
��KQ�����c��]�#�&��Il�\ ���ab������p�����썜Ü�BT,�4�� i���B"q&$ơ2 �2��HS��o~���z��z1��W�荰�֌4��`�y����t���+f.�~ρֽ?"�k�1H�Cq������q�=YjnSK�=9F�㎉X2
:v�(�x�iȌ�;���ΤMB��0k�|{��(��-A*��ܹaȅ�E<�� �����b���~�c�d�_.��tQ�	��U|�e�Ðe|�ylj`�S ��H�	�-Ǐ��)�6��}�L�N�)���mt��*aAP��(��sE�.�QS��m�]3V��!Io��~G+,�y��T-�����a�x����w�1Sh����v���6�q���׈I�~�6�N�<�mKf�W�[#5�	���J薘`q&@��isp�%W��?Mz�"\߅ǐ��������۫�����_݃O��A�=�8,�,�>R�'�$7R{a��#�SÓ�2��m�p��9_�*{�t.���vE�PVd�%�?(+��D4QRV���e;C�� j^��<��*��x!�8pX~$�y�XK�Ca�:���F��}4W<Fblʩ�u`��6������NB�q9	�j9s��@o��L-�{
���l�b��K���>�2Y�yD����qV�9���c8���Qs�D��hLt�<aq���0�fv�K�{%1U(O������б8�F�kz��;�H�J�TX�e)Q)x�,qE�<�����̒i�l�0֯�0�����.���Tʉ
�����𑳰߰���u���a���ѦPr�̾n��o?�I��� U�lI,�t���\u�m8���1�r��̮B	2��rR6B7��Q�������{�ۯ/�(�u\��\�����4�*M6��(�"Xr��u��1@fç܀��y�8l���,n�U��T�Y�HJ,)�w�Ie��ft
?�P2��0�O��&��S���)�:m[�����=�&�z�TӐ�_B �r�Ģ��S�Ю�+7�[�ᔓ���C����7Pg����&+_x���	��`l�2�T��0X	��rK�2<8����W���'7@��,�=ߓ0��_@�i��f�3[��q�R�_�#���z���[ߌ��"��Z��\K��e�Qs�Ua��a$ɧ��Y6P���Uۀ�,��C�; ]�j,E�O�!S]+B����1��_��E���F1Jn����F���Sy�Sǎ� �5-�(���i��
��f�N9Jw�c����CGLG�n����W%1�"˴z� �ӗ����!,}("�"qMv?�u��P�Jܔ�&Y�.RQE [�Im�F.q�X����<#�����G��'�1�J�T�'�妆p�;�p�1����UF\�)Ɩ7��7b��a���0�PE�43�|��!o�*��e4�������a�=PH�:@�!�_���ʫ�[�y��)�^[^v����&iZ��%�T��(Wc�3;�Aя�1چ�K�`@]�~��iP`�/5�Pq]�S�'��G�N����W�Jꪥ靌��G���[~���?���3�e���mT������d+�&&9Cd�&����ܭ�����!����o������,2��`��iZ	f���9Wi��%9��~��_�EU�e�%mB��}��?9i�Ͽªą�N����j�ap4E"�,t��`�/�䳇�ic+({�M���b�Hش8�-���dd�IL�֪z\T�4��o��������a�ᆊ[���2�ފ"�H�iőE�7	��7�9�R��V�4�?j�a�kS����14H�[p}�:d�?�'?�+������:eɾ�<IO�j�f���_�lF,�IB��k$i\k��˯��y�>�n|�Պx�n�BtO��+ K����&�G�v�fcG����X��4[�ߘ=���\�����E�2np%-��z���rو�^m}nw���� ��Ð:ݴ��`�l��>O,�	�;���I
�x��vx�U٨"_M��yղt˸[��Tǵ2���~��50�3�^�Ԑ"�Ꮠ@6�uGu8��jng��Ƕ�"Z��a��0�bzU�#+�j�P�/iKc��+��#3���=r���s�
C���l˫�D+�|H1�[�����n���Gc���W9��1�V=�u�\W�h�]��n
��P�\��X��/}�����C���Iw�!�C؄�%/��NƆ�ȑ�Q����+���!�ǿ��[����a4-[8��ї\��<�#珘4����0��Z�.�d�2����F��a������.?�/=Oe�0 �yp�G��8�`I��ۣW�mC��r�/n�Wf+��x
�?gMX��A��+�r���sD�p�:�Q&�9CSp�v��4�� �M#w����WV��/��6z���7O�Ƙ��ڭa�}����<�_�aD�ZG��-�v�����f6��o���ϱ�+`�]�d�Z&�n<�2)�^��*Q�&NB���H]���O��VǼ�Kqǯ^�ާO�'�j����/_����<M�`�(i��cH�о䳨A{0fh���?k�>z��)s~�V��4X���p^)�
�9E�����1�����ֽ{�Mm��}MҢnG��&Q�t��X
l�� ƥa8�٩m�H��6����Ŧ��Dyh��R�D=t[2���QU�s[r�{�8U�+��@��媅����A��4����C�Ƚ��%�S�*Q�A����
�����'x��Yx����l{�9=&�� �l��{k���Dmߣd���웴�iKF��n5lT�w�s(���헷�c����ᣦ̽�m�����M6V��i�BP�����;�G������o��x$wi$��ÃκL��>e���,9�⍕�t�yʓ�G���-˔�J+�����r5~�ԣ�α��� K�jx&s3�+Q	�a�Vj�$��S���;��:<Ɋ�����}�ހ��	������ݐ��M�jn���H��՚QW��,����z'5Pn�TO\�;J4��ka��n֜}���5U�W�}�7�]8]eK\�z���a�(�勧}�ҋ/X��P���#'Ϲ�-�����DÐ-3f|&4K�Ϸ��Ƨk^�|�����X��r��ϛ�a�Ð�;��Q�Tqf	�o� ���v�� Ҝ��O�W��7?^�,��5ٕ����H�u��Đ��7������rr{&I�QW/�}\���s���Ƀ$S���-�TrT���
!��(7�R�6t�>�SKf⅗�/��Z�Y��0"2*aek��{��Y3Q���C�J�b��!�S1S������\y����ڔc��0����`�.�*ӸBHè-|�ՋG���b٪�z�soCS�Y�q�z���o�3�^,au��Qml�y��t�Xh{����T,9Q��]�J���t²ZLՠ�i+:�BT����f�/�_�G�2KpP�c�	���G�1z����W	�����Z���ۊ~}���.�N��2��9��ٚ� �S�D�V�!�C3`�[ѱ�!^�g6�!��5a�|�x+np��#�$�d_�P���OB�3f���a���V���=ޤ(�O�Z��T���e"DI'B]�#��e�؈����B�Th�a���������/���� l
�����ceR�Ls�!��-"]���et��	����Q~�Y������j��: 5CH>Bq�
dGa˓W�*�/D�� �H�N�JRړ�=����3�l	2��!j�D��8�op��*�@���FM��ن?�t9�"˸(�}|��L
�|c�Ks���g�B�ϑ�.׸-�V&x��R�hO���,���2s�'+/����:�Z<�&����K��,)S��GU��l��Tl��<�F~��#�ڧd.�1NL���������SK�3���F���c8吽���"<Q�Z��
����Pf!RnqoCT�X��/gl'{ �����w����q�������1&�b(~�,��Pq~{sk
gz>JhTkE�4���V\�	��1��E� ꔃP#q��b���Y��9��Q�x��Ͽ�^�Ǥ�VL�~�b�I�<�%�����^à��*�(q���,���닆a�3q�atw6��Z&.�[�a)/�O�Ic�W_��OE��`4���g�aPK��t��R���Mq�|3�j��{y����?�+w/�/<�/���g>{�Vӱ$�y���J
 j���Kzs�҇0�y8f�upS]QD5�	�m	�!ق�y��D����Q�����fb���qD��Đ�+���(K�Ͳ8�[:硗LG���
�g  XՈ���0V��M��6b�ڒ|��ÈҒ ꑇN�:���"\5c����2�l8i�\�@ΦӢqFؘ�0sҍ8l��(���?%�Z��� �� S-g�<�n�kR+,*��N	G��1���Y��[��G���	�(R*�H�cW[����\5����W�u`ظk���?ǠS`v�m��HO�H|��4�H�����������:� Kⅻ����g��=��q�� _R6:�Ӗ
9X)�G�Dߋo��c |�D0�����	o�R��*�l�a�ݎ>���TʄdV4hiA*Q��s�+]�i���!��E��B l8���{�42Ӭ����+P�P�b>c�Sº��wPnB~u[})�z&�&��CD�Y�&X����ۯ��?�í+c���@$��ċ(�:�PP���~Ç�:��#�Uݱ>�ê� b}��x�����"nC�e��<^h80�[�����2�ǜ�c�)�O��f�N5B.NŬB4,'e���	�N���X�kx�����H��ٽa�Rs�]f���!Z�:��8�'U��y#q�vXF'�_<
�ǝ���<����OJfˠ�L!W��W56t�C�,�����[���V�|4�q�3�D&�Ze�N�@JREt�����+����2#'\��:�uA�\[��:��/���}�u\q�B`�����#N��&_�Nu�rQ���0����h��C�dJ������e�L��1p?�,�Ejy?R���pH�����G�B��C�1PV�Rg�$�D�uC�-I��-����&�Xq�CGM��`[BI��j�ֆ�	ʨ�c��1�t��8f� ��BK�p��zI���L����s�V�~��<|��}���ʴl�'$�����Q��/���c��*��	��6`�'�b���QX������_��i+���y�>�Px8�>��C���5hU��T�@L�    IDATv��/j[�|YÐ�'ӗR�ݍx�q���#���n�t��?�I�R�%�w���Y���л��KY5v�cm�|2�n��ضy�{�o�-�6@e��j��*܌�n�p�@�Iy5�F��җ�q�&���b�������y�NZ����M�v�N���d�@�i1ތ�����(5"��r���I+�a�6��W*ɺa�_
������ �,�"85]��)4�
"����YxLwiINQ�!�6�e��uQ���f���f��yU��'���
b��oy�3�j��+<�I�#�DS�uh�-ø����9y��m�I#�$�$�gV�#P��6j-]䤂����#���k:�.қ����0�ڽ��7kD��8M���1��*E�|~���.I�uN�q5���eW���Dl*�(-�2[�wcU�2�l;KXI�H�6f*��\�L鴃b!�T�VDg�b�Ȏ4K�)x�D�7 y�������G��v^A���0SҊ�����Q���l����Ɗ͒����7���8a�x��?z�Isi�aHqse�9�/]I��V/�aK�wQv}�p�TZ��n�Uf��e����7��s)�M^�@�	U+\���0ĿDj��xϗ)-x�Z�a�@x�Iƚ�����2%"|#�J�*��jh*9qY�����%�({�+.SC(�)�B"��i������^]�2T�`"���҆�D_����0�4%�,J�}��P����/H��F������E��l���\*�o\�p�=�1����Dn`+* �x%�)���[�JV��(���I-#�c�z�W-%��7�+aS�J@��@�`�l�/��YJ\���c�8�Ed�iY�XM�1����lPF�hq]�G7
�!��s�َ��[P�'�<d3�_c��-��n�3��=��T]VAɲ��	˟���YK6��G(�x��j�RN��H��*�P��(��0V���٣��{�����"�3,)����Q��R�,d�Q�U�M+Q+Hq	�j�t�|p�4t�!�����K�-���*�)T�.%���ϝ<��|��z�ghJc]QI2�(�6��&�@,+��Mtۅ��W'7�"6a�)�*'o����s�PQ����w��~.{8�c�ՠt�(OxL���*I���>��-9���B��)U򲖮g�c��0��<��6 uڮ�|�����yLɖᯠ<]�Cn %���{�*�bY����IOD*'5�J����I�9�O���I
���~�����8�I�TU�A�'��.zn����JA��Ϲ���8�5uSI>p_�]NI�ZA�c2:E���U6��A��[11q'��/:|�ra��Y�}YT���vF	;�dُ�eΐ�0�ސLSe�[�S�>�T�J�/���=��ۃ.��$TJ�"P8Q-���"5�u2�(�p]��Д˫�C�k��#�
!��Qln�ϕ8 �R���U�r�I}c)���u't��l�5!���GVg�Z:V�_DZK����;#W�s�0*
קw��`%
�+wI�It�p�M��JjE'�	p�����P��KlYS�_��JO�PjY�đ!��,�[U�7׀�AI1Ű^P�l��Q��N#�z�����qJ���W|��A�("��bI�%���dm���TTjB�Y��aC`��pR5ꁺEX��M�$E������VXB�a�{�Fs���	���<)���q_Z��Q�b�,-M��*�JY�dYF^N��ٍ�A�.��r	�Cɍ&ľ��d�#>������_B�LŇC-.�������+�oǥ� ��j���-t���lM5�%5��$��D�v)�3�BP'�7cl+�<�n I�%�r�H��������D�c!�J�c��X� D���*�8��\��ݺ�Cڑ!N�4:o�/b��*E�y(�s�i*GH�����|^Z	ZA<�DV+N�K�	�S\��+�2]�d��=w�l��x^#,ǂg����&�i��\��|N
�b���t�A)�jH-V�|G�%a��'�����Z:h��fb(���$r6+��0@���s#hl����,XF���Q���"��(A�oy���k{��C��*}S��ɤ��,&�erZ;B���6C3#)b"�M9�BH�g�34�]��r*�R2m��!� ��u�䉬�,j���؉T@6A.�T��G(����t��ư#zL�y�"�� n䢙���� �T-rVHY)��y���#��p�ɕD����p�+8_ �+�'*[�Ԭ1|��,Sl'R<;L��������\��Y(�Bx�S�\�衐;��P,Y����0ڷp�2k�!koE���L`*3-�F�F9����7���	U�#d�.̭nIT!&#���pɱ)�<ܮʺi�2Bu�٢���"���	�R)�~lp	P,�^��Z�\>&�
q����p#���b�ơ�eSY���c��)4E1�t�B�P��R7�Ur��*�&هm[s�4�L#Dѣa8r8��Ӏjzٲ���PE"�#�@���K�BB}i�E�?�&���P�&�ؕ�X�p�W��P7 ���F������&��0��'aӨ��oF��	���i�:��YzU��CN�#t���e��\C���
��ѳX�M�Ig�d��r&2`���.�ha��e갵"
�m��nظU��u���T�[���5Ǉ����a�a���(����1�����Q<�L�Z���zҠl�% a�C�ə�B�sa��<�xՖ���|��W�P(QۡNr(�����\tѣ�^H�r��l]�X[_�2����پ���|*:B���b�Qx"��͓��B�ۄ���ǡ�Bm�Z�������+��ߗ��G(4n·���y��?�U.oP3��zϬ^O�@��p��4��طe�ې��r���W=�[��;��ף�Cg�|�x�w�A��M]R.z�쁗�[����c�늌��J���{���O�0�����*ui�������L�]Y���]�RN�����s͠���c��zⵕ���ǀ��q��A��^��	��� �WF��0��1x`?4or��k�fK[K��/ۣ�ve(��1M;i��h흮�
��*�4�f��_@��Ƀ:�_o�<�V�
|��s��n�� �Y�a�]t�i�k�:|��'0�4�[?��}7\�����!���%Nxc}�B�湗�i<�*�IT�KRjVa�bȡ}1qTo��%��Qk��o�����⋿���	=�6�TzX{�!�p�/q�Q�b�y=�֫e��� �����;؝��h0P�\��ȕ!"jϬ��pr������G3�E��
Qӧ9�����{�O1�GCq�`/�=Ė���l�r˳���p���!p��/oA���e���^�V"����Si�k�1�i��3NڳRs;�:I��ت�Oվ�����}�&e"�o�ms��+n~~�%�Aˮ=/<�1~���y�yx�X��x�ݷ�ǣ�OŲe/���`�Kw����7�?��&�u�,�Q�A�.�uK03���������O���4�P�fk��z�zv��o�}�æ='?�� �&���&�C���ptg�x����p�����b՛y���ߠ��P�!ym���zbA�"M덫���s0e΋�|�m�+��߽Z��F��� ��|�࡬G��s����Q_���?���A)@�J�>[�T�!�7c��Y�}�y�hm[;@Lڃ��a�a(JQ<>����5�,7c`�z\x� �h��t�B���ۀ)�5�t0k�Op弋���>��~�Щ�߼?�w��7�ޔHےK��-f��t�s�˿�՛�j$��������]0��>�A�k?l+z�ׄ*�N�����o��Go�����ƕW��{�1v�i�h�8��#q�{bܔ���v(P��C��o���������0�(����t���Ȕ�a��`d��Kđ}�a⸓1z�C8��� �ࣿz
MZ/�4�L��'��ϋ��{��#��R���Y�w����� U�EDε�+��b���G��`����� <����۶YI���Y�ڔJ�*�GCC�p�)��ē:�򫟄�aXv=����N�|����Y+p�Q��ck�v�68���#�����^�S�d4~��!X�6��~�
�N7ԊDX���Ȱ
�n�)͍ͮ�p�1�����p�#(:�6�[ؿ�<_�z�s8x�!��I��}�r�y�x���b��0tԷ1�ʟ�SO��'�b�5� �=K����8��#pѕ�0LQ8����4�SZAHIM�oވ>=:b¨��r�
�6T&���ߏ��Fc��?}���3�����em �~7�$̜r/>3{!��yW��,Æ�!#����c4ߵ`�ɗ���n=���>r��)s�i�a(�E����I����3~	��	��Maܘ�8��G����M�*�0컇�G�,��	L��,<�Л����ix�mx`��~��V��-�p�����5�g/�OwGFKJ2͊��`�-s��T��{�`�E=1}��0;tG��ѷC��c��ᓟD���q�=qͬп�>�1���ﮧp�ȓ1lگ��O��N��u7��:[7�ǹ������a3�v_�Q;�Twdc�8� ��G@=ִ-�qż�q�-´I�`�m�����̪�Z����93��PFA�!16�r��(j�I~#�Ad�� )6�WQA�A��$�2 خb	2���9gN��f�ooa�k�y<O���o�o���U�������ˮ�h�_��폂�C���hށUs/������� ,�#P�H"Ef�^R�j��|�;��,
=4�_'�|��lF5��&^��lĶ5�u�ނYS���;_⩗_�-�]���X���֡.�桤���؉��(�ɜ1���h㞧6�t�f��D�T�7�@�9b*sp߄JQ����s���*6�F$�Y�%[8nZ��8	���7O{��è���
\��Ӟƙ��E��;`���?�d465`�X���Wo�)d���Ty�H����$R�Ԝ<�&����8��/ ��|��qr�1�:|!�pg$lb!���fa�Ⱦ��ۘ��i4
:uA}���i����w�+Y5��T���dT&$;I�q��ۋ/����w�植�N��l��]9�3z�聑����{@m��~��x�=��e/B���j�6�\$����/C	���5@���WS�:�.+M�.��^��/���kZ�9�ǅ��":�U�:�L��7���=�`~'��v���D�;�9�~֯q]���C aǝl�R�c �,����&�M�g�'�OC�)1�@N�[��_����_�� ���8n�Gu������/�@���]w\�ʝ��-@^PCYɚ��G,�h[��A�h�b������?���x�<J��F�����>5�t&o7�P,��%e"VW�ӎ;'��S�s�lM��w߆�`j9��4qF��(������a��g~->(V
�W���슛H��P:�+�Ӊ��M=I�yU�����il7"!�\t�! Yc`��j|�����'�_|�vN�]���rQTt$_�ݏ��~�Aꯨ>���d{�
�
EE��A�� %>oBN���\��t����2�G�>��O?a�?I�L�`%�����X��Zl���d�p'��D��g$-��u[�O�.֌PN������V��c��C�0���=sU)Ȑ�=��a#�#��S7�7Z�P��H.o����Ò0R-h'�nG�D
��|dH�D�3
�$d��*�����,�]e���P�ށi���g"9~�$�k�!H��$� O�Y��h���:k2�0-)�x��.|2R��P��Ɍ�K�$�3$�C�ɢHc�g/�t$`D���#�!��`�a�`F"[63�8`��z:Ú(�t>Ӏ�hJ�hױ�Ob-[��Z\͖���,�WXۢ��j@E'������I,����S�1�%f�4$�..�O� KBʰ�H�Y��:dL��.)YZ������=A�I��_h����Q$�Is�n�M���1H���a�SU0�Լ�?�d�ivj�z���_VGtU�\�J8Sj�;
�J�+����룣��b�ϝ���$��}�D"P�xV�	^�t�NӤ_J�K�=�ᙓ.1��~��č��L�#E�J�%�_P\�I�E�uN�3`mr�9V��S��G �hD�~^i�����iK�(E\�J|�t��n=��A�Fe�!�q�Rw�J1D�#{�l�4���N��7��*�ihhDT5� �GR�<$�s�1�p�Ej��bP��$b!��4!�#��ޑ���Sy�&��V~��AR��X:}!�u/DP�{���1�5����o����͒2T��Fm!��4L�:�&�i@*�+t)H1UN	�)�����P;:'Ľ��� �cW4fd�dd.���E�r���
� ���A��X�6��,�6Gy"�VEgԃ�y�Ds-l"f�izNw(�����<�"��$�!��7�0�X���Cد ������)��Mք���@���}P5���BGSFB�{o4e迉��f|��+p��/�q�o���q@�X�xŐ!��~��u���<ڣ&b>K�M�r�B�I2����&Rk�L�KuDVO%qŁx�|�D���PvҁBH�KLx�� ���[f�F�IO h5��s�t����"<j6����oݠ
�C9��~�<xD�<��A����뽨�	(��P�l&Q�y=��z�A�
�����T>�z<*)�O�r��i� �
���#1�I�>��4�KV-wׂ���]�8��/�:�;_Bp>��f`��AX����hx���EZɛ�"�[�E��ۣ- a;�G���+��I�?�I�a,���&�@��rX|:�:7㍹� f=��`n$�H�o����Ť��Fd@m��Jq�)��QKF�ʢ-�w�s/n�!�(��D�R��jT���J���Sg<�rIz󎞡��AHw�^�g#�+�e��&�q?�W�+1֔��E�7�c2��G�n�@a�
}t�/q7L����B��F����z�|�r��@��:�o*���/�Y��v�/�NG��)���v�N��=Q:�UR�%oefP�Ϡ�ڃWg�dvv�}#�-qc9�<�n��K�N���'��[�#����x��;Pc�:͊
_��M/a�ߖ��i1��j���9�����<�j�1�aĔ#��d��1�Ɣ�]�{&_rݐ���1���l�]��j�=����G
���$��AnN�H"�I�����������V�G�hE�\(�&�i�Y�G��Q����
ӟ� w���Q��4m/e�\��#�nDAf'�?8�l����+�-"F➠6W���Px�(��	;��,(�R>z?ϣ��qB5bϣ��ֲ槫Q�z)T���\2��E�m�SN��~���Dq�	�OX�z���l/�^�Ѳ`��K�J��,��~脻l�a����]���*d��i�J�Sȓh��2v�0�ټW}�{@"#�%T���$��΁T����v3)�������8��(�[[!��2��jtqvc��I�̯�'Jw[���d�Fb2J)�.��ec��� ��c8v�M�����yXWI��9zқ����j�3��l�db�Q�~�M�DW���^�}&,D����L<�����y3'^:|蠊{�%+F�������`��#���?�\�d�t�eu�[
|��1����^5���9��AWE"o4�A�:�R�T\� }�Z7�=�nԨG0��x�i @d#���$�G�N9v3
t"Z���=q`� �m��N]q^RC��G���Ǣ�	�!-�p�U���*Hd��<B�6ȨLGF;�{�il_�?P�Z��G
�b���)
t+-T=�b6�|��a1���,���<y��g�gM�lXt�ڃ��c���y�bh�����2���
6��Q����C�l��b�s  �IDATFِͪL�9̫�O����nGn��ۓ,��	c���+� �H�=�N�)G I�*�]�(���3]�`q�a�|,-C3�_a��ɀ���d .}��%�qR��ИHs
H���=��-_����j'^6��)9����<N�x�]�tw�����齿b��_Q��4���i��B$'i��k�][��̀e�^��L-DѠv�ek<}�*���0��gM��"�砆�p��qC��5���Ὕ�C�C�TB^sg��BQ������nA��5�[u/?�{��*�s=��B�"���9���$ʮ��
���l}�ށ:�I9��*�àݤ�M��J�Ŵ����x�̀�`6{�7L�������$��h2&���;����|��)9���^,A�S����a����"D�8��]�]/-㬈��4HE5��KW�b[&��(�q�5�����7,F��6Iw1-D[�.?Ʒ�h�y3�\6|h�k���ax4C%Z1u�N��o.it�g Ό�ͯ�n�}�Y�����N3f݋�Y��F���rc3�=J:����W;!)繴��+ܹ P�u\�#�k�l��x�-�U��l�d�c&��/N�	���-U������/�~�0.����EF��`(٘���<��l1F.ZP��*�~���HN��^��=�P(���pn��FL�2ŕ�d J�:i�#�X2$��ګ�������ߑ���c<�h�ء����m��
�8�:/t��n�+��v`�Q��g��(<:T����.��nhsH'���Q7s f_�d��^툤�+��jyj͕�o����i �đkVc��[������N�8}N;����"5�n��TTn�r5MX����@���c�:�^AM̮�0���[B�(Ix�����a5p�̌�2p����ɇ����ݜ60��1"���.��	}&>�_� 4��<]�	��e�fN���磋W�:����b��9=e�m�l�@P���IL����"���M�~�Hv�p�6�{/��LI�SX�2"8��<u��q��Q鈔,x@|^̊~���M��l�#Ϩ��{ou=F���ɓ�3�N�͚�A�f�uL��fl۾�5�L�.���aPZ*�ἴA���D�{A���%a�?�]lM�㟞t��#77Eg���`��񮖊�j��c,A��H7@���U~ �.�X0{��MW�Y	Sr�H��/	������p����QQ0i h��a�z�(N����F����E^$��:{i�h���PF�낳�ގ�0Zȭ�}o*g*��pD~b�a4�Q��>2�� US1f�H�:�'�3ҀM�O�6_T��j!
.��ǟ���m��6E�Dɉ����.�,�� d�a���M��B�F����9�AD�~�-��il�1��[�j��`��`*]�{�c�����h�oo�2��0�g�E-p-\�l��3�5�Ԡ��y>x��H}�(��"���3j����>�OйK�)��2"]ݼ;V- �Q��������Da~G��I9��Dݣ��Z�;�N��af����
���^����yX'��݌\���a�vL�q��ĉpꩽВLs5����4m**+w����^� �/��O�+uk!��%�'�*hH��->Z�J1�~�<����0��н�C��8�&��Q݀&L� �|u���LZ�G	���[ܶT�@G��3'�f��A�������1d���:f1��B� �"[%4�jc�H)�$2v�8���EB��x�ILA�C��+��o+�[#���m��~��ܾ��& J�R!?JXr����Q� f��#�[�`��k`�<ͮ�1����(YM�:��D�8F7�pN<�R���ɓ��˯��Ћ!��oJP���#��ʫ�z�5�����a!�ɼ~��_���|���WCs��~����׎'ۉ�1na܈�P�[���,��g�{�Z$-���j*�-�د�x`L˼{n�p��?���hђ��f�;u�b�!�!���t�N.�D��# 9̚Gmwj_s���W��p4��+��ހʏ6��:���D�@e�4f�1y9y��Q	9e��~�.|qT.k@�N�f4�"X�|����KɃ�^��8��g0:-��[K�si�L#�"��O�N�{�Yl7�<���?�v�r�(:�/�\�L�EMTQy���� 4�]i�(�L7 d7a���hx�9 ���W��W%̝>EyH;Ҏ��Ҙ~�T&���A��:f�+��˹/��5r'�����W��X��RR!`G�<<��~#�^u`������J��=��腨��9�XA�H�
zE	zBUO:k�<%w)PGn���72�US'����4�15ۑ�݁�_�q�m��|�C3|Mq�hV0�ɷ�)
����t?�$�I��a6\qxyi���T�aI�B��V-��ћ�h�4�4An�`����[;���)��ၥϠNꈌ�"��1m���w�*h+A8�#�bQ<INQ^�c#�qXB��d�64�4+�;*�D�ބ���F��iX�j�<,{�%Ȏ���g\
�[�~hQ0����b�i�6\�+y^nⲼ7Q-Ւa$�Ϟ��`����2��G��^�Z�0�����|��xR\�	�G�ܗ�Ӄ!"[p�A@��Y�rXݝ���P�8|�ǥ�uC'gBH!c+h��o6�l,[� �a�*�Ĕ�� �i*�*n��%ua�rFES�=̀^�j��'�x��_��_DpT ���3о+V��5��Ѣ��&+H�M�ׂ|}2�Z�Ȫ���b�7��N�L`!��Q��Lq�T�z9?B�j�?%cd$ah��Fg��h't҅�#�|4�R�\�LT��V��X[>�c�wЁ�K�K���Xt�臱G��L9��vQ�d��K`[����e9�V�!PR:쾴9DWd��Aq�����?V����n�nD�҆�X�h�Y_��Dn�%aD�C�0!�e'Y��[{o�%u!yo��\U�M#�To���A�b@�؃�����SKӬp"�k>m�6�H4�aPe�1�d�Z-n|�``�;:Fż,W��`��~��A<]�%�"�AH#nA�@?Y�Z\�S]�j` !��Y�7+chrr��Tj����ԓ|?���N����?��X0s�Q\��ɒ�	w,9cԃ�E���Jf�u=�bN�Ĭޔ�w��kx�"3/$��QUQ�1B�0�ڨ'��[m����%�B�ӄ��BS�x+�Ӊ̎��6��@wJ{Ncm�Hg�P뷇���!��OT@ɿ��,�X��HT�z��Ԃ�0�p� �C���1lu�Y��LC#V<j���%X��� �hT�1�n��qPA&4oBG�_��'<'�nu�j�n-8©F�6�R��:� w�V����P�v2L�B�Qj��Ϸ�4�F��ϙ���4�=;p�����9u����kR:J�!i�� ��y4�ď3� VR&W+��(7\)
⤢a^����
�=�Xa�@�"�m���q��հ:�Emb�ԋ!��R���0�.tq!�(�%�����ꋄ�th�@q^�$��MBK7C�P�/�+��?2a�
2@�.�uT2E�)��OZ�:�G"�h���O�.���,���	K��Q���I�Ȯ�߲A��NG�zo;��G#)E����� 	��j$b����"Ø;鬃�9�[�������s���!%^|"��>Z+�)�oA�����`0h�T�����+����l"S[����'�ev!OR��R��v��]ð�f���ԗ�!g�2�K܂�[�̟H[lK��k$���'霐�[Nz�.2qR'N��ĔBT|^�]Ng؁�0b��]�k��\��Y��(��@1�"�3�9�KA"���Y|>������F{�Ჟ+��ԃ�S,_>vJ�x���P{ �(6���H6��Ȥ{&�Q������;MX���g�|����[{�o�1�_�X��7�|���	r�׎)���G]R�GG���������X��"��@�K%=�MkIЬ"j
����}I�p$��=)}�v�|��7D��,�a����baL�����a���� E)����4�:+�I{����"n���g�Qk	�.�a�U7p�K�C�Ik�R6E�����D�d}��m���]����6h��io�)���AȖ�%�������:́h�[<��j�	[1�8���G�~�u��r@Ø����aCG�_���Upu�!�^7���&:>F@yT�8$�I���k?%@p�t���J��>���fh9[�E'� ��Uu8���p��I��Y��ɓ1��
�Ket�# �����1����Ҙ�S{��h����ѓ����θ��*B���+���D�{\�s��Һ�b^��E�Y* V�<cέR�<��dd,q9�I�ǘ���縮Q��������m����_��;������>x���_NsD�ḧhɧ��>��J�O<x�Fh��l����8���{�Et]W>�l�d�Q'��*�5ɤ��q'�0�w�ޱj��W�8�T��'a�R��;/���^�2�(��<�k�C���IP��C��q��a���85�����"[��������K;��Uv��=���Ϸ���_A��Y�耴�-��{03���8tȈl\�ڗ�;�zϞ�[2FWJ�e+u��訩�X��X��c��9cq�#Ѐt0(4�dI����:��a�u�i�C���2i=S>hH������믽�s�����G��T�u��*6�ߺh�/��gg4�j'�B�#� ʝ2�ʁ3���am�/���)SK��A�*�x�����������Vm��9�8�	��oWvq6֦5�/\�(RJ%�|����3h`tB��?�cٲe/�'��;w.B����ß������y��WJ?���Ej0�I_S��MCˆ����i��O<�L�/oQ�J��}���A%�Z��6������-����X���������yc����غm�i�T���%%W����c,_�ڱ�I�I#��+���?[�ֆQ^^�aƲ{R�K��۟�����ͩ�xm|e��\��ҷiVF�����]�x�0���RD�����0p������4���P<�h���'g��TTT������+��vdn�F�?��ڴƊ+��u���{6�yqq���Z�p�����k�0 �[RR�'��v��몪��2�O��hV��k+u]���a,)...�ƽ�o��*]-//�4�KZ�[%%%gfcs֭[W�u����cS4�Z�bŊe����p=�����ٸ���x�4�K[ƛ%%%����ُ���FO���n���0�b�0��������QB�eY"�YUU�@+��m�x�0�?�������o�ˆa��*�|cp�
\�	>?�F�=��ƮX��)]���c�_�|��0�m�16�������SQQ1����V�h4�+k�+W��K&���ceqq1-��s��kM�����8뮽�ھ�ؘ�k׎������0ލF�YɈܬ�]���0/..��{�O>י�yN+�������llNEE�����٭�h4zz6�v�Y]�/����=1p�@N_���˖-��,�W�b��|^66���bRee�V��v4=#k���뗴�Os0z(>��a����(�5��nݺ��n�z�g�e�UZZ���k�u]��3�@ �Ԁ?����(//�4��Z%�KJJ~��7f�ڵӪ���t�]����...�2���c�d���"]]�n��[�n��%kt]�x��?<=`��+~4�1�Y�Z峢�bzee�M�0�\��:g`nI����bN_��p�1�5M��CT���������0V��P�yXƲe˞�,����&�V����5�\��^Ɇn۴i��P(�m�T*�NYYY6�յ�a��y^E!��篺��~4�Ix¶��4z�r������|޲e˖�Y��DjL����Ҭ����� �G��~���k��u(>���X�d�R ��(�|��ʊalذa��͛gAZ:�&5�#G��e�ʲe�^�m�"�G\�OF���� V�\9'�J]o���ܹm�ϖ��e�Y�f͠>�����;��pgհa�f�0V�XQ��'I4k�����,���+'fk�o�sXy����Ζe��i�i���e��nݺm����ܹ�g�i�h��b�f�QG՘��w��A����$Ɇa4���U�=b�Z��6���Q%�H~��8�<�!ڃ�����92f,    IEND�B`�PK   ���X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   �z�X�H2�    /   images/9865acd8-fab0-4625-b565-b7238dff6b6e.png��PNG

   IHDR   d   d   p�T   	pHYs  ��  ��F��   tEXtSoftware www.inkscape.org��<  �IDATx��]	tTU���{���JB��H����(���Ӷs�>��n������\����e���rfZg����E�dI �'��m��VD�@UI}��V�{�����WUWd��+l�zsWaV�A�&���Ա�6K�
��9͆�k����qmE�M�th&:�d����d|Q=+E�i��Y�ڈh�ɘ7�����ja���:�|kq�C�)ƫ�'�m�aӅ�)ߋ��:o#��yI�!EA9�j�#��q[�l������
��"	a2n]�?�^�n���B�%�t�*��+������������x��y�=�)ܟ�PxP��e�.�1]��C�,��
���}�TG�/'r=7r���`ܷ������K��*��y�n�IWJ��͚�S��+>��ȪK�h�I�����]�?\�a��!��',�o"|Kѱ�tԻ������VN���K�����ɭ�Q���b��Ah
z`�y���/����#H���)���(pI��ֈt4R���w ��9�ĄL�����T����{!G�?NY�B���F�:�� <N�j���z���?�Zy��Ɓ�t$�&��#�m@�'��5蹝Ɉv����F���^�mm"����-}ʉfiw[�<:u��Y<�o2��s��z�$���~z�g��[M��Asȃ�wL�?m��cs���ikA� iFi���<��!�ɸ(� ~?�s�&mW�Y���o����K���Ha��� ��������Ćj;�\� ��L��e�n鷧z����?��*�����W͍_$ᶄ�u��zY����N�T�\��L_�O/+؟����N��:Rɠ�p.Z)M*짛y�N��ˬ��yKq��݈ʖH&^��3(�Zb��he)�y�/��T����e����������R�Ť9cf�������%ס����fp߃SZ��i�4nxz�
���i�y�k�"���乼`?HFmK6�>O�e���6��d�Ҍ���F�8�(GV��*��7��t!��C �����9)�vJ7�*�HO�a�����rf��b,� �|��Q����ｺh/��4�
6.�9�����6�rW�#fi�����2�?v���/(.��!�UH/W���R�O�e�d:�_\>�'�����Lu~��^a�N}a9bZ6f��?dbK�AM=�{d�pPDJ�sg�w_ɘ 4#Щ��zx�C��U�F�!������
э���8���_�NZ�ϐ��ᛂ�9B�m�m~Y�TU���v6��>�Pu\�޼�6� �}�PU���t.�����ၞ�PR}��T����ܺpס��R�K�:��	WΤ�����@u��LM�Ec�cG�!l�W�#?�{d���r���`�ۺ���.�-�Ң�N(�yE-�<i���;�N�a��)ퟆ�ݔN�r�T8n�T�%�%{���HK��/�Ŝ!��v?U�%踓��gJ���i ��8?�k�IB�h�ӹ��[��2d�T&�4�L�4�!�2����N}9M��Dx"�5�Q���x��:b'��r5��&>߱̦��:��eCȥ2�h�}Y���:L�e�0b��,� �fN�5dӿ�
�%ſ,�X�l��4�J֑��Œ6���[+7ȶ��7vL�f$?��!�֮�*>�Yykȡ/�?\&R�)1}���[�leۂ4��A�iË[Γv�����i�i����?��h�J�t<6Q�����`��?p�e��4G��f�&_��4�41D�w��Ji~�c��=ұ�p~2n[	ˊ8]��j`Y6��t�if��߯=DQs!*[S�W�]��ǵĿ[;�7�`�VB�Z&��T�i���(s7N3L��3��~ |t�'g���Zu����hx�+s�_����@
�)ܕ���t<��|RY�,��*XJ���J<r�&Mn(�^��k��<E^�#�fҦ�.����.ʫ�c��͔Q��+���DD�2aٰ�(�z�ue �%�R���`�Q��l�ƨ�s�_ˇ���l���(KO�����o������8Ni�G/����$��3�C8��6"��x��B��nhC���)c$UD�ᰦ�+*�gm����Z��O�Ɗv�df��\��@u}�F�����1*[�$�@M��������6��$�0n�d�Q9�4Z�J����z���BT�~ؿ�.��Z�8,����%d�F����
���dȼi%���i�Hc����ý;�]���<v���5��_!;����j��)��0淌I�^���;�G�Bv��d��fz	j�ڰ���� ��KŊm�1�h0���G�����������L�cR�r��_����ٟ�1� ��'�����P���l��MuL3��٩TY%2*1o�JKF�WÁ�Fh�χˆe����_�A9����H�%m��s�L�f�n�H��d0��
6�^C���|���Mxh���k��}t���QMu�t�F���6T��O��b�v�aG��3�Ѐ�u͘l:�RY���E�ihF��fLQ��� t|��uM()� +��Ɂ�rQ\�G���:9vUC�?�MP� ��6e�u����ADZ#T4P���*��&�����q����p8Ι/�x4.��Ҧ\<|ކ�Ӳk^�(ʖ闣����
ß%�`��L]�K죇�^�^����^�R�$P�A����MA��G��IY�:��_ʵ��+,�/�B��J��u�p `�`�}ƊU.t��&9\~g��JAsY&��z+Wq[ZZ�眂�;�il�e�M���;�Φ>�_3z���-��Cٻ���A-I�|u~/v�"�����tMA@�����&�˷����q-���w`��J��p�6���6�k�a�d��<%l���`&�s ��SH�U��V�{n<�{������DHNv����}�eH�A�&"�������^�D�F����ț��ɉ+J�:��F8��:�߉�]�R�B��	���F��e��c�smM%�9����%��3���5����!��5��9�w�	BB"�\��=�>C���:��ν��i��P�TV�b}��-Ӵ�ZK�!}!�S�0�=�s����w����m�9B����8I�.:��$!�%	Bb�!��g	a��";��(�iB�QK�4!�xӒ>OHXK�'���0�)���ē��B����O3�5.^�����~C#V��!�%L
?ĊU�+B��XV�~ұ��O��P(6?���aD}I,~��_��08���o	�D�?�m�ؓ�~KC�"���5yz�ׄ�7p�t�҇��5!�h+��%� Q�*	B"`-���*&��3x&%<�|���-��>�J�x<���93]	B��sm��t����s��� �0�H9��+A�	������N;�5�x�1�� �.]w`�f��CA�?�؉���4�q���	�e���������Gu"�ȑ#���E�F������$w"$���?k�W ��#%)/�k�(�J$��5��?B�ǃ�Ay�m�v���B�	z?C����~����x������cw�o+&�X�0�^�����k����I&X��|�?w��֫��b�!.'(*�6�A��!5o��zz�:�+\8+�=�C�mIƍ�����>$Ɛ $Ɛ $Ɛ $Ɛ $Ɛ $Ɛ $Ɛ $� ���n�Qb8i���tu"�\�f�g�y�B�Pyw�.61�e����28����jD��sd��I8�^$��M�y#_�>�7Eh��׼s%oYj�����P�WR8\	������Z,A"#���ҳp:�lGE��T�� ���d˲<L2���y3IEqe�̅�>�,�媼�0n����7�O�y�B�m)�p�0�Y:UrG��l_�k�C&�m�j���x�o�,$O��n��4�N���M�q��m����T�U�M���o������^���^~wa�
2��xf�r\S��'�JR�Ť1��ee�͙�Y�ÛF�Lyp�|��g��^�mQ�@�y��k�ދX��?B�U������� �17���]����p��v�s2TM�"P���|��y__�>�^�%Bخy��W�}���[���[�]d��7t���������>���K��[jw{�h�Y�
ϐQ1O�Q���v���l��d����>D�Ͽ�o�?!B�:�!My�4c�5���٧Y~��*�N�ϸw��L�0����fd>�w��T%2tem�~U��틧f�*�q���>J��HM��c<�^72������h'�W�+贻��~Q��[������nSx_\A�֒RRM�-"������}ءq�![<:=��������"�8v���Ɉf�x�8.��8/����~1�������"�"&d�b�ff�����;F
iŧ��?g����*��Ɛ�^~�#P���{`0wp4��KՈ�HF��QI
��;)-��Ϭ���
]u�$�r9�\(LJ&��6zY1$��H=usű�r:(�p�֦b*�B������Cض�c'�8�e�2%TP��ߝ����Ք���t��L=��2��\!?�xj��#6�T���'�вa)ڶ�Z�'�m�ʗȎ/J�8;��o�x�T�Z���'u��l���T�mJ���'�I�����q��a��ߨ�G;�)��%�'�PB0�08g*1���O�=���ɮ�.�"Ye���Xv]iIt򓟙�0��>|��Kh�"����Ua�3�Y6��.��B	�-��1�ӪB��O�dI�v��G������$�o��:���2a�<4y� �ڷخ�� �HJ�p���ROv���,Ƀ����aZv�Ŷ�����Sr���N�<��Gvn����ww����#,�$�c�5f�	���}#����	�Tג�񹨕�.>��1M����K['�^x(f^\>/n=N��$9�<:��NI�»1����CXOo:���pݬ3�h�IN�c��|k�
~��<w�2*X�z~N͒�%~n��"Ҟc_Ǣ|%_S�_�q��|@0����g�h��&m�/���;Ғ5�*:��U�)AG����x��9���82;��^L��Q�X�nc^�b�����݅�2�*,3Y�����n��4b�
wf]�����)d�&K�3A�g��l�����XP\�qa^�ՙ^?;|�8������d����h�},���ɸs��thn�k��̺�<ɉ��|,�f��l��_��K�D��x�    IEND�B`�PK   }�X��$W� >� /   images/a4664b0c-b4f7-4551-a44a-c7f07c5873cd.png�USL��{��Ipww��q׍���	����]�����]���9�T}]��gf�u�Z�J���! A@@|��W�����_ ����X���߁� ���:���L�C%�����Qs�:3;��^�fkjNkr����!~C�L���#����"�o����8G���#2��0g�\�.j(C�ZxT_����w5��}�U���z~�p��-nn������������g��H"y�?�L5�� ��O���:fQ��=3B4�c�`�"l��B)������A�r��w���#�?��#�?��#��Q������
<��N(w� I�r��WT]�ܳ�h��=v�4������
�� �FM(b��5ӎ�Z��:a{�9Z4���8��Y��O�7�xY#S�HC'Tu�h�����)8ݿ:��C~��r�K��4��u��B�w�m����V��B����y}��gG�{�R
���f��O�<2�����{N�i�����T$O��D��Z� ���������<���:� 1� u.�=�w*�k�*��u����	}�Pm�\=֒Fk��3��$��z�]E��u��%�*�ųG�X��b�y!����L�� �����$�.mf~���-2f~�o��%���_:�BW�!��	%Q��En�&�]p����zy_�L��/m�����J������tl,{a�2՘A��z�jx<���|�z�N�]4���mZ���s4b����%��LJ�]Z���֗K�1�/\a�K¦U�A���Ѷ��:�]U��k�����dv����G���b�G��ޢ^(� �2]9ݭ���Z�Go-�;,�$�O�������됛���� �ڤ��	�:�e$g]>���?��rL�(C�;3:�	utm��qO�:+��D]���J���ls��CȲ����3���Q����%/������n�=���V���S��f��4�֫�j��x�4m�NK`�]���m����6��0�m,��c���=�������ڝ�Q�(?{���T2���E�U�2:��$L��B%��V�4L���}w���O����>�Z�Tf+u�Ŋ?cUK��"9�����;Ñ�e�o(�$��-�ΟA��d5�	��&cS�dao�4+�{h�9�c��9&:]��Q64m=5,�`?D_}1�t�a��Hg^��h��;9�H!W����&����;($�j�Y	�^�v�v��1�=��fib��[.�aHy�)-��Fm�8
�P�y�q����X��N��A7Mh,���S��������������w� �&i�4�f�O�G��~���<EV��9/���	xo|�W�=���s{S��o�e�a��Ӌ��im�����J�=«5$�ԜJol}�������\~Ȭ?�8�E�R�G���iψrZiF� IG���+~���h;��i�^P�օ�5p�L������gZ�Q�����T�+�.�+]AY��|�4j�����MB�DƘ �Z��0���5���F�t��)�H�-�=Ty��jD��a.����C?�]�x�Tx� �	����;R�}Y�<2�1�!q�\�+�~� ���A�?��L��e�l�:�k���ǂr�7����h͑L&I:X�~lOzUug�]5b��Ɂ|Sl��ʃ
�=����worn�q��h)�s��o<��\2Y.',���	ٌ ��~t��#�jg.[�b�Y�/J~�OǙd��~��g��H��¥g�.z�:\1L.�׻��s��~ȳ��)�칁������ۓ���]��ߖ��F+�û+���/�V�n�����bLl�ubW������ ��0i��f��c���,. 5��tU�x�@)�T���v�i�R���t�c���!��{]�,�:2�|�
�I�MKn����09�w��7;���O�/��.�RQ'�Y���%��gF��d��_��k=wi��F��i�)�g�l�KQǅ��\&�l���������Sʠ��y��zYjF"�l�JQF������T�TБƠ�~���h��O?$8�ѷz����a��PUJb�������}1�me�4xfw�S����^��m| ���kW��S��s��s�l ����W)�7�8➪ۢ��έ�[�; ��!h��}�>�7^��[�=��P�b�M4�m�	�G����M��M���@��~�bZ�&3ڬ5I��u��q������N��]�,ڃ��X3 ��9��:�ܳR�9b����G�$�\�#K"e�ÕI͈��f�/X�2������\Î�l���ޕ��Bt�����n�¥z'��� ��~#�YC���1�	�L#A���ݻ���|�KK,�D�[Da���V�����
��M�j��Z��(D?�DDKZ���E����D��!�9ʚ7��'��=16�V�Y3������������J�� �G.B$B&1���j.'�رm^S�4�x��ھ��-֖o���=����"AusPNؿ^�$�Nϒʁ����f OW�
ǐo���8h+y,�wѤ�'z )ކ�?"����b�!��;FS��d;?��1V���9M���?�}���;c��(�xը�Bj#hA�K�iJ<<���`�k�J��=����N$��! �iE�R�@���R:eO�&c\uF\�T�=�@�_�k�Rbo�N�Zõ��	y�_o37�7Y�� �D����ew��_as�6L��uE"1�2�����1����ս��Ș���+m8̹��&��]i��e�4���G,v� �K."�P�ȟ������c7�9!���<p8��$��&Ձ���Gl�[�l2	�?��+Ual�LW������q�\����?�;�J�YS(o����S��m��r�uI��ʰy����Zְk̦|r�?�f���BE���/�ƛh���/��޵��Ӝ�5s3��y�m?|�;���/o���o-ܰ�E)���:fbUj����
VK�,݌J	����FPٰ��^�.]�<�2��Ж��wa*��� �<����K��EZ��#.S�uR�n][�T�I�%'gg��0cH!����|4����0zNw�ې���N�� %2�k��k2�

��9F��A����I�>��N�|CbH�cф�^���i��ˇ%u��o�:�7�L
@
�	��G	z8��
�@�l���'��l��^��Q넠��L]�^��u�	Hۖ�dDQ�MKY�^ต=� �����$�^���|T�Q�0���9i�C�I['C��l�l�#S�_)/A|�snx���<������=G�q��\���B�z� a�,���'Q���2������D�ƙ�}\ô�������)��YJ?�5���Y�"E�E�(OOO0�'�#?0V4�!Pb�_I)4������>����A?�y�&�b�6���@6ᰉ܇@���m�����Ai�Zy��N_A,?,ϡ�g]��H��?Ux��c2�&pro����#W:��y��Ij�ʵ���y���N
�âD����`1`��+��#k���6���Y02C��u����׶�z�ԯ4��ڙL���/�����/%c�Ǵ��x&���"SL���/�Yr���~�3Q1�0�9�B�~()�+.��%$g�l6}�4��:ZG��+�����1��'�ݥC�	(N+�9�m2%G��t�;�n-uʒ��� ���z�j����z��s�����6��]P�YTd��4�>oϹ{���-�;1]�I���H��y�"ܥ��{s�)p.А����ٗ��}rzo��y�7E	 ����]�!���z�8���*�*��������g�.�	eI�j�W�a��2��߂�ըe��;R-��@-�f$���-��YEAJ�(��N�c��++�����.�l�,
�V��7[�MH�C��+K_�}��O�B�A��H��`��G�'I����		��鍖5"v���J�x{K�_&7�g��>�1RFg�)ߔC�!�;�s����2���l��U�0`;���ԅ���(V2���U�-��C�%M�G�M����*=y&���\Ҭw��"���e7|��r^u��kNY9)�b�Eb�.!��Hڊd��v�Ҹ�'��c[���Q�Rv4���%p|;q�
G_�B5,{�M�����QN0����T�T8ұ���_ɔQ ���j8���=\��h���\�U�$?��w튡Z��Ϊ[a�Pw�:�!s�UQ�{F�	;��3)��t@�j㣦�H��d�����7����҃��xo�� ���4?����d|E��y8q�aec���Q�8���#8`���<p�u�7�?]�
FN��x�T
����2��j�nK�P��1e��&�k��:Qֿhޏ!���J�_�%V7�ҩ� ���GjU+8]�"ް^�v�2u�6��:� ��/�b��i%Rs�r}U�f�9EK��oW�1�F�d%��]��JsGf��:�t��N�?9��͙-k~�$7myb�à���
�%��:��s,]����ܬ��SG�2xo�W�n�ا�r:f�_����E�~>@u��@�ы{2]�>��*�YJ�2��#���!�E�F��(F`39d��7��+��n�[�L����@��K))�% Ob�A��ҡ� ?���/��� k�%}.T��!}�:T#bz2� $��j�i|�o���m}N�r���y���)
)9p�A��SMU��Y�Z���e�H���o�
�s���4��B��Q�k��Y��щ�g�6�C��	�@꧖<�5E��5��$!�:�+Vm�O�B��lx����Ɠ`�̟L��tA�S7�O��n�c��?����d3�tY����V!���m(K-�!C�Ei��C��*t�21oa�;].Vp�T@B��:����S��&{jPЯo�S�_$5|<�����JV�޻�:�eG^I���(��l���!�)<���g�<�ŃX�K��o�D
T#�$��f|rFѿJ�������WW�Ph��È���@�*ys!cG���OxH��`�Obb#A���5%��ތ�~���d���x����_��;���Y��W��ע���,U�jgj}��6[��_�cӌ⽝��ؑu�B>�x���Z��A@+��
�P��;}��@�}^�e|m��"��_X���Ҡ!����y_�X�_}L�K�`ZA
�Y��i7�H�y��[��O�YtC���z���SC������ff����-���^S?���i��^��n	�Vs�LQo��ý�ڏ��H�&3�C�JI�t�k|��ȿ��i�
������*�>1��^�Eu�%ԭ�oHO���jJ����/�I�tr�R�s�(E=�l���<��";z�;V~Q��~��tL����-�r'��ܯp7H��$Rqr#�ª� f��w��Q$�cN"X'����O��k��`M�=%���_�:���/�(�hTx�Ѧv?�4�O�`�,ꨟ��YΛy��j�p5�E7�����Cw+���A��"!9F4̨|���y��ܣ��`����F���q)m	)Q���Yb'd/���\���9�sj���5��:ZU�B�~4z�M$?��ᴚ�R��/"|�ft1nҏ�i��&C�<���ۊ���"
�����b@��0�?ٺï0[==�����!V��(��\����ڡ	k�����MM���e�.����c1��7v�ʯ�(/	��$R5����N&�L���L@3v�p�WI�����T�,o\��!����29��[:Y��WqΪ����[�L�En0�Ag�Sy֨�]�����M<=��KyLe�I��H_�DJ�ԑ��0y- C�v���p�i�I𭬪�%5V$Yo�[��2ɦy�����?�I�T��p
~�G�n�)yP��7��D���Mb��LH��;��y#�ޟI� %�o�u�/���� |a|�QgE�LcC��jU���Q��X�o��D��,����-�g1i��x$2�B(a^p����n��N�@��i��Ο��-�e��y#�sd�O���L��H���h*�gߛ�i��Q.�p`y5t��vn�T?��0m�_7P�姢�-�r����G��,O���ܸ�h;��|���]ḯ`m�T����CNw���}�`��>O`�Xe��򑯒=ħFI�]/`;����l�y�{?� �����%!|��n���yIۣ��[�a.&CFO֌�%�#�H�V�P��p��R��m�`���>���H���f��������A�>�������C��5�3p�g몍^���W��7��o��Iu�?����{"�XJi!�'J
?S<=d�A�D�8�R�``�m�ǃ'�~[�q�p�\�n�"z�%����%66�!�Y_����BL��Aow�F��N
@c"�X��V'�A�J�Sz���G�6�Q��zqy�sIP"a�e�+	�v����Eq����Qo���noƄ�fxz\���~.�W�k�a�;|�x8�%-Q0W.e
u%ȕ;�\!��3c)�͜�����ZuW��Ue��=h�=Ts*mfMB�o�g��]�+����h�*X�E%�k�5HF$LN\�L#��(*���j\���?�pJ�O�i���lCo��o��ۻA�#���a����b���DR�B��y�#ф/&�L�T�W`Rnͬ���q����▄+�p{4hc}NC,��tN'6:�a|��D��hA1m�V�2e��"��9
��˗�ePכo\�G�$5�"��"q��`<k�z�-�-]n*���-oȬ���|����V��b�.����.�XT~��t�x�nY��I�c�.����/����-�W����V4�rt1cV�>ǋ�M	�T�!��)Ǖre�L�Irh(��@/��n6�g��^�u2Ut%q�I�Pp ��
yǴ���+�g}�1��{����{�g�(;Q�(Eq�#?���gY��p��DC9�C_�R�?��5�@ho��FtoHN۸�S���$�����c��9�[7C	��z�ֈj�����0-�:r'���guڡ�B�u1�I����H�-�ְS�_;�M-Yv�[C�V3�`M탅���yz}���@@�/��3�����f��{h�h��Ә�V��rS���^(�(�k�:�m�����,�+��	�*W���dt���(�X������f}M����}5]�_F�D������)'lIF���I�?����82����Y�i%}�J�\�q���I_ĝ���K*eL�̑!⊻���>9�§�)NSz{�U�	�g���	Qm�0ŵ�Ƃ[�/9�F����0���H��]E�
M7�t��c�;sdJ"����%lTb��+D�>^��	����Qk��V��׎�Yg�)T�9�L\�O0r���ڨz�p���5��C�"%[�V�
�ܷ
5졭����Ԟg+
ʨP &E����;�aq����g���ֻ:O�w#�|S����+_��.R���jW�� Qgֲe�B�P�:���|���q�T�C���KIц=������ͫ�n�n��snFy���Y,ٹ�F>�S4J����P۰d]�_�@?����6:i�M畓�ⵉa��m{�6UӶ�����@U^��#�$�
���;8ւ:��.�j�t���2��tޣ9yNg����I�c�ײGꆝ�N��PV�ajbO<�.�f���jSl��ͫŮ%�Y:Rb �n� ��o=�Y�*��	��9�����
�$�#����I��L��2�r*��0+��/����
p��9��mkU���-�&��Vj%K����,6��pteZ�����	f�`��2�=a^bw��A`N�-�YXZc�ăԭ%hT��F\J�\H�Of:���z��L�����h��rݽ���~~V���q��o����Vd6%�>���Y�
J�%MHd�-W+]Mp��r���l�*�J��Z�)Vw����x�C3��>d��1-��%K��jYčTLz
�o�@B�]���xC;�W=��@���f��[��O83�ר�.�B�p*"a�FL�O�EȰ5}��ui�e��K��=F�Af��LB"R7�����/j�����9�oRb�*˲0�1�)��e-n�g�S`��k���u0e!�z��ϛWC�h:KN�Ή������刾U7����m��X�+�����No�k��jy���wԼ�El2E��?�'zn�>��[|]������1u?��u31�<�t���1l`r���ӧw�C���Ũ���}�Β
�zY�~�l� �Ç=O=�]���*x����[D�e]O�/�|+�z��fΞ8Cd�l)�ei�Z4�|*1fҗ�eà	�%L�K*;�y0� a[9�-Sig�O�������/�mv"�������,�"�S����|�i�*��wG����[�" ��mŭ^�l���ֺ����f�����۩A��{j	+px���@�@9���#s�0���G �y3�|j�ũ���]K7�#�0����#��N��~}�)_����ʿ�WQ�Ds��Xvz��ʍL7MZR��Lz�|v�Z�S�nP�ojBVpL[nɁk8$e�@'��H����cט��"v��ރE�ȯ�M/6�4D-����ܙ������)I$b��A�3��V7��\?Ⱦ�XR�����I��p����?M1��?��Qk��cE0���J?�>*�X��6���<%��]\��6��'�&�%�UJ,:�f�:��h1^�fʸ��:�aR&�t"��e�]�3�CaU��F�s ����c�44b�72*���pnn�jk;i�P&ze�Ex(q`5R��V�>HaB��<B�;��2��P�?ԋ�[�U:�w��ם�+݌�<=���8�M'[ˑm�:,0�}�H�&�к����ٺ�F�{yA�,ge͌1�*ΐ�+�-���G63qK��Ao�+�E0	�Q�\�9Vf�"e�K�����I�hH�&���S��Ū��*ok?z�
<?4��� 5SX�S�Ȕ�����}M����$z�<�B��������ά8��UFy��b8�WcwtC�T@�ʫY��t�q��tkc-k�r����p�k��x'<������h���e>V�Oi��,A|u�#�8g=i0ۇ�r'���"t�� OG����� � �#6!�tǞ���6���qɝ']N!�L����I|C��F�w�{x+��1%���;jl�f~�����=��v��F���J�Ԛ̮��f�qNCG^�G+x�8��f��vgO���/E:7�ф����7g]�%���oYگG�8�R4�"븲�@����2(>��_��J�5Ya�3㠰N��^O[xl�WLh$�3��a~��
	��U�ɗ?��dQJ���U6>L���E��m�_��8..���bP�m�!?�_��O�#�8�/k���9�YT��S�C�����؉�S4G`W�R�>G$xiy:��B"�-Ǣ,ŝ���H3�0�2l��$�����ѡ��I�,7�bz�Q�Ob�!��,�93����"��S{��B�z���Fuay�w���u4E��(�a/XK�A�8��IG:�S>\#�O�Ϊ �.��(|b�W������
�����(*�U�Y�v-�n��r�����]W�oX]}���<�胈��S?X��,��P�����:��m��z��H��p�a���8�_�pF���+EK�}� �M�iFP��I��i�{��A�p7��~m�����Q#�;�T|��Ѽ���s'݄��8��&{3����Z����1H���[�Z��#U��ћq�F	�I]��H$i/�&�N�|���t��"[�䰑��ъ_�TC,$Ӵ��^f�I��Ծ�l�/���A�퐂�$`����4��4Ll��f�� �k. j:��4;��T�}]�
ߕ��G�e���ie��j��!��K�߸L/�h�we*E��*��,Ddf����U���.e�!	�ыR��<����i'�u4����~��j�9sۥ�΂�~pf����L\�-��8�Fc�^@���w�O���,{�DD���[Y����вb�]�V�egp�|���l*�\���ʌ�e]�
�W0�7�a���|���Q\;�R�&#�)�0�:a1�v�`Ԕh蝨��5+`�)8��$^� K.��+����'Y�7�掦���qRz�nCe����H���L��|��[�w�UK��\��N�̢"�e>`�c�`g4��G�?G��UլeE�vŐ��Gg�Qk�R0�$����iY�?I�ZN;�������8$���4�V(T�z��Z�_�R��'�C�1<Ye"�SmjX@��`!�0eNF�f�H���j�t�oY�^���as��)!�UV�� mI1�~��0>:��BzvQ�Gs�V����� �C��w*K-����fd@,5M.k���*��*ɴx$+P��AosE1o�����2��B�`�J/��
~����'����$�	^�Rl���%Ǐ^���i���e�������ԝ�7�}�g�!
�����tu�Wh�XS H5&����af��K��Ө�5��k"������tZe#<v昕N��Ɍ�Q�z>�Ӎ�(`��eτKqQ���;���-	.��֕XWo�ѕY��g�������JNi�Y��&����!s8dX�Ēu87Dp����q�7q��f_�Q�c�)#������ 1 Q�>��O�\u�ڜ܆+����O^c�V�$�,���߈�"��M�D�D���u+�Fa�6�1���A���������B)�8+��;����[�3j�
�\�ߕ�����;2�)nT�Z�HM�Թ�T�T��Jud!�ϋN�A�C3��_�y��C)��?����_�PjOP�Ե��<��[�ד���:
ӏ�2��;R�VB�E��E[�H���Y|�h�U�[�n]�4U��7�d���BQ+,5("ue��)=�ct�ٸ~�É���H�����aӹ��9��9��H~ڎM��8k#yC�eQΚ�������-������=j1����r_��{�3BZ�:�P٭H&�a��G %�w	����,Vm3���PZ��*ܮ'��%�ڿlu̧>H�죀�S<V��V�|��1&���Jݗ�I�(	����G���"#�U�00f�A�)�^1/��Te@�c�g�k�m�Ŀ��g���8{��P�p2�gx�4׫m��Jܔ��u�����/jܔ����.,�AF�*o��N..ycf�5r�M���p���=L����g�)!	޺
�������6���7z�:�_��JH�Z�1`�m텊Jb ���������SgZ������mb.��R���l���KCV�gf1[:��]:�gy��s��1 x+�p6�S�8���"7�����g%��F����4��R:vL�]��\�F1���K ],����|���̙hv�Nv_\�n���'�NϏ8ơQ~vZ�����5�@�B���K/v���v�bekD�٣l}#8�9���X�Y^#�>�����D�9��:�"��ǐr���B�m��n��c��])-� �"�\(O]���BA<�u\e����.3a�/'d�5�L�sKy�B�ģh�=4$�Vօ���	�$�<ip��nG����Usz���6���?6���E����-��L�"d#�.,i���v /�ɔ�o��*�լ,K�e2�N�TeЫ 1kB�%e�ʚ�#���H/'�`���2�n���DH�K^��kیdX��rr[}l��E�ECr�0=A>n�r�بtzږfPII�}X�v�~U�x��}i�Ғ3�,_r��g�|����[\�u᫑�z)���5����ȵ���y߰��#�Phj+Ƌ����G@�OW��^�uy�|E����Iۓnr΄�6��}9�>����:��N��/��++�;Nx���9��x�8$�,��+�������A1a��e�b�@ �ڙ�?T��#�E(o�H�l+b�n���|���t�� S�d�V�0��=4̣�r�r�Rfܡ+�@v�Շux긋��w������a�}��P�&d_�
9=�s�؈���35޺�ߵh��
��� 4+֌ݿel�z��."�y�����w��G�%�,?0VfqLڅ���էep�����pmy���y��9�z�D�1}�6V����
�kA<��VD�|JN�.#;ΕqƬueM������0x(Ӵ$��c���B�������qSu��?�2W��ॢ���'!�^����B��k�;���zۖŬ���U
s8F���Kh����c���/Kn=��N�#e�S{�%��{a=N,jG��]�`���\Y1��~T��.4�}'�T <]W����~B\t�3�1%�kԃ��1Z�l1]^��isu1N�+"-���q���} 24.�~��KE�X���8d�Ӭo	����fn��� �;��;z �+�P�kf>9:J��ɔI�
/fV�Q�7m���٘,�,3-�XlL�@��b�+���S�y7��1w�#�H����Ex��	���ƴZQ����saM���v)��ەɪ!�Yo/L �3W3T�3��dL[��p/�Ec��&s:��T�N�R��k�ҁ�P�PX��)��F��$Qs$�-H��~R�&�����3�Թ�N��F����J�g��M.��פ�[�hː�K����Zr`����YJp8�T���ʰz(�����XO�tcg�d�JD�9t2�ͽ���<u�`eq1��fKO�aV�^��1qT:�|R�i��ު���d9��Yaȑ3ۚX�-�<#%z0�t��#�(��h_���"���㯼cO��z�ߢ�	�C��f�d�gC�No��+�oNd����tt�B�qՊ���-	V�B+a�?J���%�HX�j�F�O�`%+�@	{J��R�D�k0�*�,�ax�ǈ�����GGIB�f��b�}��,�!����)ΎQ"^��Vp����zzFI��a�f�aT�`���w�A�H�H'"�X��j��/-y;��8q�(H�j]ت�F��t�@�eg;��	��n:���B�B��f�?<N&��{&:��;�g��ͨ�_��tq����ʡ�{:H�~�x��5�{uo�^��W5]ZE���2�/���;�?��p�J�݉�9�d{=��@n�mC�6a�g`�9Z����x��I��ß�Z$P�Y�Vt����KsN���A4�w9��am����tzx�yer��c!�7�m_��3�3���6L�I��T��k�:C'	�N���g��ہ���,·���%�f�̂��צ܃�g!�y�H+U�)�p~�)�Iw�=D�q����)��D��$W%��w����������4�`����	/5��e	W����H+#���E_�wf5����+�-f1�>ncI_O=P���F�����6��F��="!&��De�(��U{ca��u!{xȭ}!�x����Jvf�|M�B���{�J�5�{�[Yjw�E�F'B��eI6Gě���i���CS���b?r��z����p�
����|Rg�8��ː7�Ub�Ù�&tо��ǂ�i��S��H�v����(�7�-v�p)bn�m���x�56iѬd�Kh��$�9�P�N�~Hx\��섑��vݒ$u��V��R���X����k}�N�HK�v9Ѿ���8vG:�":���]���̴�J4n6�'*׍�\zF�R9!%�G\YGq9Q��Zt��:����v`]�Au5:�#�ԇ��G�F���ܨ��ǯ���k�M#�j_t�d��k�2n�C8Z�2��qr�`�l�e���Kq���<��ĴT��{O59�m\�����;�$f뭴9�=���Y${�O��F �����x6�6��F7/2�DK��ҀU�֭�*����O�0��[#����	��J��g[K����Rg�>+�����=�4/;�~��Zp���k��8���e�`B)��3�	��	�rW����hs~���s':�/o�2��}
�� hL[�},���|����aeZ�j��+��(�^�Zi�e.9��aT�[��vo=[U������_mv���mɫM1`Epأ��:�W�WL�l����ݴ'J�_�I�X��a!C�}V�{6��	a�;��e](���[_���#�x�ݫ�'⭧/�;��Ƌj�	n�_����F"��8+N0�����y�x�׽�(�����1R�
�~���r�?��� �δ=i�55��W�^��;b-_�gp�{�DWW�W[�bm.��E�s.O�|Y���$Z���r��d9i#$^�9�<^�T���7�?�{h;¤�����Ym�?��ċ,�:$�3���Xg�5���5�O�Z�2����dҔ3�ei��;��*
��h�*ȥũu��Z�:�UVOuѰ���r�>� �=a�bPH�-H��f����~��<!=��&�����p���ib���^?�(����l��z��t��7=d��|�(߼���?�	�C*^��\����������,k��c�	��[:,E�jW�2�kx�7[��U�� ��]�R�i�C�q8w�E�]��	s����C����݂���u(ea����� �pP���e��7_Wۏ��ŭ��ROYZ��uD�{I>ڣi�Ƨ�f���R~�a�4��i��D9�7c����Rj���B������'Y�
>�T
9�,I��f`/�|�V ����׻��q�e�c�n��VM_�e�m=����g��h����%�^�1�k�D��r�S�]Ys�3M�G2�������ZLe�9�[�eekd���~9��Ϙ�u��z��n_6RU���|,|��?�溏�4���WCy�g]un�A�Г�Nȿ����&1�H�|��,J�e��W	�g\�=�D4(�����DLZ��Qf�P��imZ�Pz	��'뼅d+W'&(絹D��4������r���@P�xY�@�Ɖ�<���7���)o*���2ў#ו�3�>(�Aζ�>
�ԏWn�[��i��.m�5r�A|I͢�� "�2�z� vt�|2���
z�z�fz9�sr�_
���<G��Q�g��!N�왆^L��6�%���r�
��暜�����2:���мY��u�j 綛BK.߾7�/�؛	�}���ftȵ��Ov�����i�!��\�<���(�/xaq`��q%>�7�i�{����N)9����>��RL��}A��͌V�E߭�
c3�{2���<;�h4�Z�㲍y��p�w�f�����Ld�"�������=���5���t/�#a�����Bۋ7 �R�g+��]�AI�����+/���) ���U`�X3l�1k|����Df㖃a�
�h�u'��%<��Ԭ#UbdjJ�X�vy���Yr׼�B	\�^b9޻<<��<D���W��k@+���H���Vɛ!�(�a�ᢜ��GB�\�O���)IF�z� ���S����a�˲�i2Rbb ��b���I��. ��fo�W�� ��_�{6��d3Ea�Cy�oM����@X1���"济���>a���/��1Y���6Z��{=g��q)�8�M'���^萳o��̈�y�e���v&�r�2������&܏�8?oz/*$7��7m�J�lbK��x�ӹ2 >,�my<1x��Ҥ;�։�=;����F7�j�8W]m\�S*�g����ͩԊb�P�W\��h6T�R�����?$�j}����;��T�N�|���^w�ʋĶ�� ���\�!���;<U5ju���*ty�)*/R��q1n�@��	˥�l�!���=��t�x�YƲV�$8c�ˁe��┗D��NZ�^[�wN���#���Z��Z��-����T��S��+\����QIf��&a�s)�[Epq`��8潝�k�5�E�ފKV�s�k��N��5�OT�����]���$���s�ƒ��|��4�L��ju�؞�r�>���>V�n7;,�[U�NK&2SdN�J�U���A3�U��)�2�4u��F�J������<����55V�I�L�� ��m�|4jg������嚴���|<�9�5#w}	�썫����4+/UgO�g�K_@;���
�%��e7v�a*J���ņ�gc\_�a>wzWhj��
b<0�u0����^V�B�Z�;��c���͓ŀ��һ�h�C�1��<�%�i���c�M��bm��pV;PaR��@�"�����Bc�ή��Fk�C_���1ϥQ
o���6@ɿ�/Wm�ݹ�+�h�'=T��gu�Z�[�#X�s��e�	��C]����4~̼�6���l�:H�L:cyVwe]���P6�P(xJ��,�L:<ͯ�N�N1ߞ�^=�=n]��~��[OT��@7��ܹ�k��b�����r}+�;������E�J(��P�޻{[��V��?!=(!c�z��T��?�ģx�H���uZ�o-�,��������G���zK�tIPj��H�B�}k�ZV��{�.z�����`"o�	-�m��*b���Px�_��&Ǉ��daJ{ɻ�ѝ��63���#��@F%�k�k��B�ͅj���ϊ �װ�X�Ϟ߂)і�n4�Z&�;�eI,'�`�o�����������Pݲ%�����X]{���Ez/�i2]�4YȔ�`q^����s��C�;݆ ��o����G/i��_����h�9I�	N�S��]��s��5��\Ȥ�u}}U�n�j�K�Ν;'�wMΞ=/gN�SM�Νmi�yO�9+�����D��N�xk1qnrZ/,�a_����,�n,���*:�\}_��?�3�ݿ��0�Z�IX��׾"������Y�({{�R���`�&�]�b}��`Y�`R����s!;ܩ�^4#�c@2k{tQc�y8��PF�K��Q�ꔮ��.g��}l�cgٳ��4������I*m_��:s|�,gKک�T ���W$겟�΀���.�\ۊ�4�9ujS3�'���s�qG��\�����+�x��L���Y�$�\����2T���yF��4aN�,�Mw��M
y�%]����툾9j���(�%�,�;wwdeuÝ=��\����[Q�"�ㅼ�����+�8"׋ O]9c�7����*�s<��H�A�L�\L�:Oƻ�R�y��-(��F~xx ��؝"��k�2fk���H��7�뚄Ɠ��ݎ6~�Gc=�n� 1�k[�q�*��O&lμg��{w�����=3`�*	n1����`B��eG�2u�2ޛ���1e㗮63����W������o���җ�RA�T�AІ:t���7����;�j�:���$���� ;f���!/�D�c]q�QvL��d�[�\�8k�Dw���N1E��ǅ�2o���äJv�l��i������O����
�2յ�J���Kk,�1��> ���$`�1V2��|�`���f�B�?8��:�2���a,�t�i�!�0w��$w�}��-���o��GR@H�SwO���n�;�\QK��5a�ם�TA(��]���B���\�XU�9���o���k	�8,ċg��H�Ν�r��$]䲶�ɒ<���ݾ7�2��/`��oo+%2鷳�U���y��G�?ڕ����#��te�º�y�Iz����&�������zmI ���ҥ���d?3�y����P&�T���Zb�kK�����G�������O?��<~墼xkJˊf�=�����kݵ��eh�R�P�0l�`ݢ�&�HŚ]MRb�	��tϻ�1��񎌏v0�,BR�x0��ͥ��K<=ӝy1��dSk��/C�����.�P��)�[-�9O�
5�eF�b�ּ���s��KZ��-f��k���zٔ�7�)�N���C)[;-[���99���*N
��2�g���P=��A���193ӺB��O,���n�H����˙Ñb���vD�zf]g�\5����@	�xk����Ң���?c�Y�{$�F7��C�("�\�ɘ�#�#<��O%<�ݕ����]mi\��xz�VY�0�b<�4����\8� 6O"n���k��>��ꮭ�p�P�p$zc�t`~i�WȲɝ�(�w��60~�~B��@Z��o�]�l:U������US���\�tng�N�����uUZ�P�� �o|�Z��iX�Q��ev<Rw�!��?���������SU����ʍ%u�C&���^=�8���c���0�H���;bf�B�m!O��]!ͧ�\�'5�㦝t����!�s��XE�fnOF���`oMqmr����i�(��2Tee�oY�c��}�JS�٢�ӾH�����
Z�l�R��$H��l"�~��y�-/�;#��@��ҙLY�� Ync���UX������L�y���I��<�J� ��M��j��ei?��g�kǲ��ȥ���D˫� Ɨ_~Uv��iH�Օ/]�O=��̦Z���Xa��K7w��D6�dt(wnސ8up���;Z�.�Ѿ|⑋�$6Z�	��W����wV�;����@>��0����Ԇ!�x��<)�|��t~M�x�M�~��dOp�?����㟽��Z���/�D��
��l���OR~x�;��^��;������9��%��$�W�����%~���Nz�R��6DL��B��p��br 3�X3�}(OQ5�^��JK��[	���$I/�h\B�[ф��Ka�B���5�k��>�#Y3N�&+�1�csE	z��%�we��� �	������l��ʹ�e�1�u̖������������$Q�e���8�K~�{�V�� r��Z&{jWBV7ຬT`l��-Q!�q?����r��)ia�B�����m%����BpvkS�$lϺ�}Anܹ�I��T�y��_Uk";8�W��@֝o��I�랆r��Z�/��G���תzC2MRd�9�	��!��'{P�\���%2,̙{F���թ�&���e�$��U)h�6�&t�������>�-ݭSz ����ݾ*�t��Z��~yM�
=�8��U����-��U(;w�������X���{�w�c쳶�ؼ��[�3�֑�Z.����r�"a9sH+�ɹX;ܫN�i�>��'�+��J=���_�'��5�99+��qa�d��i^=M�Ŗf;���cMŗI�>"{�"��>r��Ҽ�Cn�le�جY�����i�J_
��}���Pc��{(��x=ơ '����!�n`�N�qM����Q-o�4�Z7cĚ�w�����E�}��T�ja���luB9{���k7�>�M���cl�~�-�.�5ަ\<FO�*����_�Ek2�AHvCMRk�n ÕB"�*��ӣ�Z*�bߥJ��V�sŧC��qo�Noh���<��y��̩�t��[s=:4f�q�`X�T4`=��g?���yN>��O�w����v�C��6�59΃�8�Փе\J]��@O'��A��n�띂1�c#E�!��i)²�1��5,�b�ubY�Ų�	�(a�X2�f�3�M^�;���w4�Qz�I1�<�&��F�lȐ�i��ӽ���Wk<�<-��UY?uV�&gXO�$i��xv8=ц$ފx=�)ƛ
@��ϽUv����W��|q�������^�]cE�jZ��X�J��4Ù!�B��!C%	�/+XO��P���Nb��%�v����t�Ib���持L-~m
�l�U�肏��̑�0j�O?����G/���|�[ߒG�"O<��6b����Y�MW~�v�� �g$[_�](\��P.���1� {*�l5��\����x%O?�4Iѕ��޷N��\�{�c���W�8��Wz�|���kOS�����~Ҫ��t����au;��	�X�J��=��Ⓩ?!�=�����r��-���>�_��_�_��ߖˏ=!�g�P���9t�>$g~q�VOB�k�n�`Oz8�t���8zj�'�P~Ͽ�<S�MO�c�&4�~OR<C��[Dm٥��I�݁v��Nή��O����nן��rxr�Z3Wŝ�$M��_��y�?���/»u떏�������������w�����Ś�yN^�.>�H�,S��8�	���ϋz�
(�3�?���
��cVa;��i]NϞ-�=�T�?��>P�i�T��4�` �i
k�-H}.~h�1�@������a��}U��=Y�v��)_8Դ��d�����MY��	U�/��*n����eY�kB�_�@VV6��ҊUX�3%��Q�̂5���`!��R�
D/g�]K{t�����cA`<��CODē� �Y���Zk�Y����ī�ݦ�}\����fC)�s��E-{TSi؀�[?����X�q�l�1�A&x���[�Z�Eza�s����W_�O�����ӥK�Ԣ⑝���5'J9hܫ\�3w~���W}uyR`;���ߔ�;�`�Lru���	
<G������!��Z���.CO�P��T@��Al�7�`�/��P�]�-Iʑ���=�wM��#��mD�>��l�:';�GX#3MRs	~�
wZW�V>�%k:zT�<s-��Z�B���������W������&a6�l��ԟayz����D'�Wo��@?>
t�F f*m�|Ci�ky$?FK�ԅR9����Y��>ݮ���Q���\P1{�ɧ�s�����?�c9>>�?��?-$g&5�_�K�g���_R�Xߐ;Ñ�w�Yd
��
ȍA�f8��H���
o����j�6������y�����1�J�H3A��jd\66�d�;�7�]kē�^�@�0�Y�	>k�0�L��o�����s�_��"o����2�#ƺ#�����B�@�{��um�8�п�ͣ0����^]�uba��zװ]3�'ć�mU��{��e���֖~����yJԓ�A�9�p	�
���3r�AQa�)��,ue�nT��ot���8�Y���n�ū�3�����x}�%(X�Ѐ��L�P��V���WP�)�L^E@��b�m�̫6�~�f0�A�ZD�ͩ���5�y��u��*�/6 ���/���ٲ���v:��{nNݷs: h�@�H��ȑ4URyj��~q���R�jF��`���v�G�D�I�@#h�n�F�t��tr���Z��O_P6,@�\�Q�o:g����[+��Q忣��ȳm�H�{0����~P��,S,�EY��T��42c�OGT1FL �K����k�c���~�˲~7x�|<p�_�@2�!a��Te�^#D��]�M�L�@��-�˖f��f�NqL��@��
��� ��!�đ-�f�#g$��Q?�gt��̹��^p5=�@���#������U�L��|��i58#%��Ȏ��a`]˨(A�9�H3��(�c	j��a���$0s�X�0���B�]�z���P�y_��z�W�e�F	:re�H�1���$��=�j�L�8��x�̜�k��=�Wd 3jTjbDa��t�e�ʅ�2c2� ��W����0g1�JX䆻��л�\?@��]̪S�PG>�Yވ~������5���Mv�ң('�������$5hI�n�/v3$)� ��]@�kE��fؚ=�4Ӷ�=|���<ţsj`1��x�k���p1F�0(݃��ՑoJ��Ē�¬81ޖm�(�X)�J1�L��:!!.|"���Ț�M�`pN��ݘ��c1v�����x-b!CcL�sh��׉15<�>����Ը�J27;Og>56�q2t����k5f�p��RA>�v_�[˲݇? Fƕz'` ܁>b���	h�  h���>�giJܐd: �w겵]c��
�i��;h�d
t�̘�V�s� 4`�V&N���5p ��P����)�������7�d`d����l����ζ<v��|��):t$4{���M� ��b'�$ I"j�o]3%��!zo���eaaA�?��p�h�I�_p�Z��,ݹ)�ʎ��y�<V 2������܌�	p��v��*���cG-^c=��u�n�*�	���$	Q<��'�hIb�߶l#@�/�GN�a�=��5!�����h༝�J��(V I&nl��������wӚ��d:)�n}�w��F��X�7��ȿ�����~����G=p�_��#4��)v�#@B�F�jA�A(�������'�o�nX�|P���	�<��&3�)}1�t�赙�g@�Xd��6�$�S���r5v5�^][�i;\��L �^� \�H!@�̢����G�Xn�Zx_c�4FP!�1	P�)7M���r�K��e�5P���
=]�i�W�ɍ5�����B-�~h#�B�����`��}*�� ��`�l�Ga���n6�m��i�Gԣ[XV�`���
��<��-�l:=�.��p�yu���iu�Z
)p���ӨBd�g�Y��^f1v������*��5AR�E�QKz}��#;zT�-�Ƿ�d�2bY�ޑ�@�!h��>C��s �9n�	D��@>�u���T�sH�a�9�����b�8C3���vr��>�*a�I��COÚ#�=u�nh2m�bKy�g��K&gڤ b!([8p���w�ܚ�p���o��@�T�]c/|��7/����$57k�Buhm���n���
�N��|��(��W�{SQG�rxs�!#�j�$E�.x�Sb��͔B��='�G�^��j*���\��7n�>���f"��g�z�q���txhY����Z3bAu)4{��P��
���읛��q�3���2G��p/_�,7�]��}3t��^� Dq@FH��P}��T{'ub�.�	�\��r�;���"���?N:a=U��'�^"C2�k�18ꚼ�q�="�U�gߨ�9M5�Ҧ�5��B�R��+�2dPýk'�m��@d?�iA��8~�0Vvc�)^Ǧ ��2�|e��X	���?���VD	�t�������*��D�x�F�6���v^aLt��RV������;��=��K���^F� ���� �蚅��M�DA��VG�eR��:��Z��btEl`�� $1��v�O�cJK�2���D�˧�Ź��H��-�^�}.�1��ؑ9��υhq\%�c�3��h���>���|%.��&���9S��'��0j,h�\40���́�f�y5��PA�.�����އ4=�SY���}Ȇ:�Z�,�k��RٓJ30�w�ng�M�j�� �/��AG�n0�pT�;�D�ϯ]�H���>��ޣ���ԧ�����M�&<����:T&K��5���ጣI���Y��g�"�33)O>�W��������6|�W7������k�Oه���T���¸P�x���q]��@,��b(o|������Iv�&�qb�peuIv6���׳��L��PK �H��ǂ����d5��b�m�; ���쬈����b�N�(H���}�`.~�I�:1��8ݍ���o^co����JybZ��O��s�`[�~����wHT�H\R>}�m\�:�>�灛�u��k��_�!t(Y�AW�#�8�̎�g8_P:Cr��1��0�z{�ժ��A|Iv��}�g
��F+�%k j����=��s ��L�=t�:P+�=�!���u)�sG����F
h�k=1;+{���1��O���cc	S�} ��(�`��WDUE\�c�'fH�aJ&�������=vg���z�X���i�A��T��0��M�b��(fh�(�c��b�Sv��/���d�ؼ��<v��10����q�NX�p~14�ٿ�Fߝ1[��:Q��{����ц�h_����z�I�v�G�+(�iH��n�'!�b꩔�,�ߗ�������q]�!*v��N%�ހr���&ەf��VǘF*�l��b�h�HSNH~z�<�vfv��j=nn���f$�K4�V�XH���˔�B�p�m�")%��Ō18�3S+@83P6:&bOțh��'=8���K���Ǳ��10A��!]��A�zwP��FM��f�s�i�dimK�'E�2��:Ri�����@Ô_=�����N��l�ާp`�Fv��M5B��t1�c�e��p�%�LvV_@,ߏ�"�˄�Ǐ�)��7���U�x����d�UÜ	%_.I���)��y�jk;��V�)mK�i���D&+@��'����I5�ȑ�QYک�zeG3�2i^@�/�]��<�620�����8R��O���!+���D�	�<����Q'��Ե*�m2���7�a�z��&8��S(!w�{W�e����Ё�@\�6�k�����T�۷���TJ�����o2�gA2��h�J׊�R��u3�s��I1�}�;����A)ȹ_�"�/]��%���y�(5��R�\��5���qbU�W�F�8f]�Z�j@'��Ee"����J��E`;��[��ޣ��rYÞ��,Ld{�S��O{6���������i� ��S�{��P�> ��S����^^� j�g�?���y����z/R����2=9��oU>��x�D{L?L��F�	���>�%�gS�>'�[,��i�LjH���e�a�'�<q����z�`YN8;��� "�B�Y���ā�Qh*F�ӻ��:Ѥ'�s�8x�w��߃^�m�(���b���3�"{��cF�K��G�ʺͷ٢2:�NL�e&�8��DbC�,�{�;P�⊂�(hP�������/�������C�V=�s��F�p7]�0�pA;	�2��gɾ�Q9y�	f��}��\���F�)�'=�֨�-FRF:y"������:�!p$˦#�4W���E�+e|rBR���f��k-dx�k�d2CSFc_NY��~�?����� .��Yb&�q�|��ЇG#Nxd"}��C�ϲk{���f�+�)���m`�� ����I�e�p��P	3T�0���w�6K���Y��i:���q˔�\s^��1��f�Z��������O�4�`Ԃ��W<:�[*�N]R]"O�V��b[�=k���G�efn�#R8G��aH��nW*rO3�b8�F�ű*�7?#���P6��I�Փc�Z[Վ,֠\�d��gҕ�f��j͌�&dT�
���힡��'D���!H�F�SD���Iz|�y��YF��R�V�O.~,-�b�x��D��w�۬�<"9�ك����;�~���efj��z��.�tzq)ۢ0��ƎT[�XU�3��	.����my�ͷ����?��>���TQ���ɓ�o��3ې�:�Fg�D�e��"������o��m���҆ E�?��pj��M9��o��SS�-�w�y� /�ڴ��^��E
�h6Ց	
˗Fy=������Ir���Q_6�7����ʮ��Ǿ���$���R�葓�ѣGc������Ϭml˿��O����ڂ�t�"c����=��2Z z������(ܛ����}�BZ\�I���5��RF��ǿ�Mk@�*ZڜU��6D_#{�(¤	���o��#0���6��T�L�3���n���l�	?�> ���LHo�*�ڋ�iW2��?7��H�4��Lٮzc�{�j�:(�&�G61&�����1�o١�Zz�BR���4�m߶l(C�A-�'����}=���y�v�j�Z��͌�^�������T�x���8�/q �����Ĥ
Ԡ-�23��6�N�@FG��7�27Z���xD#{��~[�^���H0� �	�]��,2R���е�L
�Qp��D���6�0��:ʣ���G6�g�/pc!�{��d��޵���>�-w�_�� /����,���(��쓢ӷ��0�y��\ۚ!t�5��@�B/޲2,�64��}�)�6RAC&�i�̪��5�,͐��Ꮻc�@6?����W�Q޹�(����N�L�]RD�& ��S�Ե�`�d�C��h� �u���
n�nĎ4Y�0G+V[ ���Z]^"��������� ;_��$���cϕ%a ֐�A`C刮���xL���N}S��H��fG4��s�l	��"r��C�K��ߖ#�e}�ȹ� ��K��ʓ@r��!��çҝ����3ױa��L�9^@bXK ��桡W�2hw�f.]��68LV K19=%w��d�A�dyvd��<��~@оC6;�.D�|��z#�".|��dYyṧ����26=+���V ��j���XT��s�5";m��,y.���ruC>�s��.�k豷���yǧ�ĩ����/s�Օر!������m�~>��e4��"Z3 h��9�uC �)X��i`�A���}����u����벬�(`�NM�������Λ�X�+^Z�IЏ�,難o�8Bn�Ш� �2�)���p&;���5�uR�K��]����E�X]�{Kw5Z�X� z�1�h���T$��;�Ps�pUoƖ.�A�uC��� 
�j���<��C7#2������:@�k���y@�X�rlL9u]�=8xֆ��q���ߪ���~��}z���Z�e�T�Y��$LU�Zss��WpݾZ�y�X{=�����Y�;4��Ĝ� �TJ� D���a6;Ф=���pP(�z�{'O��U>�C��.8o�+��^��D�c�d�7s�%n�#Ƀ�#
zn|D�G�'27R�Q�Ǩi]��"D��vH'e��-.�0p%�c��������֎T4�Z(���d塇���� �e{m��W�Ɛ%�Jq�a>�7us6x��7 �"�O˂�3���$�'����M�y�����	�_�ߔ^e�Ղ��QIזd�����������,:���)����6��ݿ�E3��-S{��j�R����u���xr K�D�g(va��b�mH��]u��ʧ5��5���!Y�75� (bDJ��� qml�&��w����f�N�8S��n^�.]V�@G���`{��內��	7u}�;���T�1��X�$�k�
*6p!˕M���jX�@�F(��/I"�ax��$ ��LD_/�7����6���7�T�1�� ��N�i���#��� ���@����xd�dypP�i�Tȗ�fQ���OɊf�̸<�r�L�s!� :��m�o�um����1�ކ��9�~�A*�+f,.�v�I�	�*��=���絣ϵ�ϡ�� %�>lȂB� ��^c�Q��k�g�2u��^�lT�/��V@������]}&���~9̽��v��� ��k W��`>�oA�=��f�6EoP�#m3�U>��siTkb��"���hI��tA�;gp�ρ�O�+�b�4�u�m=�����z��\�r�0�8#~�g[����UeЂ=��{���`"�#��u��
�ܝ�H��F�rf|�f.�n[�H�>-]��[�Yp�t�i��,�S�$���F���nǉ��A4H��T�R)�����4\L��~����o����}�Ư�ί�6����@i����C�GH�fd@C�P��5`���ufALP��)��˥�Z����.��<��P�̸Ԅq_'��!ч��+���щ*P�04�;��dV��|IP0��ձcG��w~��4�w �Q#�	d�ƭl!/�Iڻ�kZ�&x�2
Q��ύ��.����w��Ր���"�f�lT��-�4��L^�~,�x2��dv� ����\)-E�f4SO��zN9����3'	ȃ#�r��P~�v��s`T������f�4J����@ S ���Q�P�:E������ۮ����Pb��K�T��$Y����7���%���q������k��	6��ߏ�~\���/3ӓT�c[�]��ջ����;�R~�AD=�xHk�j��W*�1=´+;��4A+��/�g�ἩI��M���to��l\�x�챜�n�1B7"��t8�3���}[G���=���8����Yg�Q=vXnܹc��zώ;&Ӻ.���X��������!M�Pq(�� �[��HV�7�7����D� '����ˆ��� oЦ7 D�~,iF�駟JD��,��-7�S�݁���Y۪�k8� 0��q�kD��@̨`S,lE9�>.�4(ܔ�������՛�_���A��h�c�	P���g�{VF��6��QG�;N[1�{vM����|���U=�"ZA$<2זTq$ ߤ<�̢����=��jK��Ɍ�?�"��w �Ny�D�^�@�k�4���G�D�}S�卣���ѩ�O���K[���ʎ�KV2O!�G�'��Yl��)�=��RR�A��g�P�d- \ɡǙvY�F2Yi��Hc��8Y��
��Ԟ��b��� �%*���+W���D}�fKyy������^�z~��][DOOO@DG�繹�i���@�:]�tqN�zkX��y仾�R�8S�=�Z鑔��J�ΫsWûU�fuG��iVZ
���'%�sd������x���9K��a�>v_Z��L��'O>rƔ5�YY�'�o���l��4�Q��Q$�ݲ�����	a���i�F�g&_Էl�5�k\� �}��d��V����$�`&��B.O�rE���V�Jj���2l�P��9=�ٙY�я~$�N�2Z��k��rO�+BMI���0��#kt6>1A�Nr�8��U$f�vr���>&�s����x�}�� � �=z�Ȓ혀��*1@/���WA��
UH���t�`F�Í�Up�x�<a����D�&9�P X5>V��|"j�c�yln�#O�O�t>�5�#[����g��
Y�͒{��&\Y�5��U=��2�65�򡻀2�������S�={��kۧb�G�]컞:�K��X�Ǡ�)P�C0�L�7���q�㣣2U.3()��܇@���-r�Q���x8����ٲZi�i_�x�,2w8e����o%�:��P��ȑc\;����g��y�U9��eFq� k�$�3�p�����q����Nz�vW�q�-a��D!�5���t&�w��H3[�ow��a1ӑ�1UL[���"��3[���%������8�B �>[��1��	�.�5J���Б}2�w%�%�ސ}S�Pa���M��'�������T�9��'҃.q�l���#$OY7���8��D=���^���ՙG��.9y�!����'����dcC?��g��N���������z�N�ȍzG��i�V���v��5f���#��ދ\I�PF֏�O�\�Mٹw[rj�\5��^FZ�Hf���H��o�Ug���7��<}�!���u��ɧ,9��=��e�#f,F���ؤ�h*�V<�4?�uH���'�"���ô�6����pd&�O�$5�I������1|�p�@Sm�r��2<�8��@H7�O��:qR^z�[t�nJ��k�;��H�:!3Hd<�j4���,�Y65��i/�Y1?kȃ�g�ئ+/2�꘤h@A$�|�"�J%cLt�1"Z�-2� -���9�{4@�:��9��/\��؜����%�����6j��^�h��8�TA��<����|)C���Q�6�����\.�w�������O>���#���ӧ�f��^{U�O��Ŭ;Y�� ;���Uo�8*��ьO��L�=���ɔ����QD(�V|��,9��)��^���		z]�u\ݽwW����:�c��3O2 �TK__`�Ғ7߿ �}.[Պaecp�NV��+7���n�f�YuҐԝ���?��.��������GׯJ�^c�C�Y�9c:f�;vrt���i��ə�=�A&�6�KM����J0$���>J�=z2R�K��!�?�-t?�P��=�o��_�����C͘����W��9���׍0���关�DAd���c���6l_�-����t�4kبud}�.˫k���`��<�0�� sa)�6���ű|f���{}+��~��y94=)�����ɲf�wn���d]�|�m�	�ia�;�������KO@>*j�����fü�fRj�;Ӏ!l��1�o^Z���TmFp�P��UiOLJ������d��=��[ӭ�K��r���C���ߢA��r����J�e:���X�]2΅��jl'����>�>bV�C��9v�!{h�D-f���G��l1/�����einX��
�=�#�ļv"�&��e�: ��!#�.����ظa��L3�u����y] '�:?�
�<9F��٦S,���*���"�zVߔ���GE�%����m�̦���8���U��w�6�h|��At�����]Y�'��V�`��!'Z!�&|��W8����\O���d�p*�nn�Ґ˦eϾR��w�����?}�|���5�l���:Z*u�A�R��o����,���4��2��G��瞓O?�$O<��<�����׍�* U�k�/_}U,��"�$�P�� ��ᑲ�8��o��P�J��tfԮi����/Ͼ�iU�e��mNm�8��V�~���{\���]Z�Ԁ���y@�3{���P~��yu���zM(WHm�� �8P}ސ!�Ԫ&��5���t*K�,RT�Ǒd�I�� �Ȑ�=a�=���1�/����FV1M�M�L���
�2d��%4�\�ۂ��5� 5�^ȧ���=���x�п��FN��.z��0��|�}Ȍ�d)/3#j����P�Kl�1�n"��hrɏ�����cjb\jM�r�,f?|�XB���Lx�Mm��JA��f,O<rJfgNK�A�`L���/�s��'~,��u�@���ŸX�(5;;۔���4�{�#+E����JS$Nw4�A�LqF���JK�x����Y��Sن�D:+E5�Ⱦ!汦���Tϖϯ^1 <3/��	y����񧟕C�������ȝ{k|M
D��3J�:|&	�E��7d��+�&�!�đ������9`RJ��xYr�;�Yu���I��%kK˲���ƺF�z��9pdpj Wsh�'�:�t`�-..���4{�@E���nvrJzV[��.�Kh�nv �e�mY1��f? �\��Df��0f�E�Z�I�j�Byl�r�Βv�-5u<ӓC]y��s���������^?wN>B���mѩ�`��|��\Ӥ4����kM�G�x t�~�T����ʟ��?�ɩy��k��k�10r�yߺ��7���4���uև�9>F�N�G'�W�`������Lk;����l�o�~W�٢^oZ��d}F9	��R�y����;3L:�9��]�J��!C�������'o�~���談�	dbzV�6+�W�K�́��ԣO�w�Cy�3r�T��3wS1�KFF4�,k�>�!܃B�(/��2�g?����mpd̘���ʒ^�=u즢�0�!QHh`N�6��I����4A�'�@"ޓ��|T;��@�`�>�Ӏ2�������%���;�������8��b�7*�9��B2�s�sƦAO����%ٿ1+�%���I����Td�RZȕʎDj($?"Uu~��^���m�	��c���b�G`�U)J��22�h&�ƿ��_IY��:$%u��d�G?���s�᧗��as���Жefj�%� �Zu�aܬ�ׄ�'��d����H�Gu9b��#/m�cz]�{@r|L�i\1Ǜ���G��Lv�mJF�¸fk������Y �4�����\�zGz�WԪ�����3i�8k���V��S ��Db�֡(��ħ�$z�~W�΀���S�;�����YHN��3s���Ƶkr��5����7�B2��:�/>/;F��9���}��7��@�Y�!A��Ȩ:T]Wu~~Q����jK�`W��G�z�����u|�& �4�LA0c�$/
h��o0���8.x���q������)���>q��i@�oY��=tP����Ҷ���f½���U� `���	���������c��6Dpp�sy~����������H�ؙG����s���v]�3�@������?��?�ɱQ���{�Z3^N0� `@uIF��oa.����e��]�+�r��)�� X,�2�G ���c��F��<<s0�������C@�g���Ɓ�g��m4�gf���>�k���%�զ~\�L�$ߍ~_��Ok@�_�2�x4��o� /<��L�G,C�6�3���ſ�`�Mu��)H���u4`lp��hېT��&�P����L��<{��'$R	��p?��-�d����F�'$��S�J���gXLk���_׭� d48	PX������T��K4.C��N"�n�%d������|���M���ʀ����E|9��_�~�{�?�\^��k�Տ�:%��׶Ը��|��F��1�r�}�}KSN�9��\�n���y���K��ӧ�3�/���� B@��<��R����렏�X�D�>�3��f��s���,��g��/_y�T#�A� ű�F�K�\���5+�b��/�+0�b�<K���6�uJB�5�o5Z��	�Hf�&���������Yk�&�`l��)Ns��xª'�]ʉGւ�� �g�rY[pő<��}�TT($�� ��=���ޣ��y9r�9rB�'ߓʶ:PI2��8�Ѩ��Y��{w�����A�>�P����hW�TA�/L�xjJ֝1i_���Vd>�9��$C��~&i� �����17�O!tsO��P��F�ԯ0𽾡5u]�gM�'30��I#�FYtQ����'��㳁(����Ac��Ē�XW���0�nq�m�g���{2l���GVAt݌��E���]`�=R{�7* �@\
�#BK	��L.-=\F�JrꑳR�t.�̀Wx��[o�VZ�:��8���L���B �1j
 �@.�_��ܾ}W<�G5=�pY̡P!�
���Y�o#�o��2�����c�k%.�ooU�#x���ek�"}�s5��H�۳s�r��A�V�e��-�л�F ޤ�F��>'\Q�w8���-�}���A��KN�����0�CJaDʘ=���%0����x���xp[��j(�J�2d�m�W
DkF3��Kd5t�_]�J�׈�U�I5��c�f���ت5像>�[2#�	3��t�ژeb)2��ɸS���I��'�>v
���O�H؈Xj �/�˹�>fO��Ò���,=˂���I���L���|H.�����f�(՟�pQꚉ�GF.g�qN�O���s/~��6�8��q�ߌ���NtT����a��B�Ҭ	�iqy[��ࢼ��yY�ܒt�,�f�n��m�Y[7�)t
^�}"�����I��� u��
�+��@�$@k���������� �-mjd�E��4��@�H�є��ߕ��Ui�k���Pd�xf8�,Fx�it5s�����?+˂f��ʜZ�QרĹ��n��@�)�P��β:�nt���M��a���h����S�F��=����`��#Z���8@�L0��-�h9��jfG��������f�������R!���Œ!D�뺱���r���)��h�� �AL�2�w�x��u��i}��<��St��k��@�W�ْ��I�Pg
�_�M�e��Je[�9s��Wq}���\ZY�t6+g{T& j�{� ��lI�c�C��E$����6	2b0��s�n�,�2CYX����E�G�(��5���F�\3���\��wޑ�~�`U@N	��@�;x��4�N�� (2̊������>��1Aƀ6���g�!���f���VBR����w����hG4�h����+��!�0&a Z5��Y/�H�_�����#�B/��Ь����@�NL����Fh�����|�Ź2:���鄦��!q�'\��b�Kc\]�v#��шS���Dԋ�-�S�agI��:*�Q��	��o�p������-[��<r��L�T�70�0D.G!�+�C�h�Y�����S&3Ao���y����y��/�Ȁ�X���R���cGV���<�����0c��dj�)�д4C���r{iC�|����Uu�;R��O3�H��2|s1���02��!�e� ��E�[��i�$ P��m*$��M���&Ȑ��� ��RF.�C��f����T��hӎ�cxY���P�2�#�`X�c%�
��VV�Y�XۻG����;>/��(pF8�M�����l��ҧ��.�A�� J����$Pێu_	J��r�h3���pu��a�U�ֿ�|Ƴst-�|e6d߳���d�����a������-:-��	��?��������J�T�|���W�^�����&%`O=��_SSD����%(�ϩ#]����[poff��w �A�<��61�}���"���W���׮����_�*&���3`�ԑu���r���v���>[4�u��k��������D�=7ְf��`���`(�(�.\��|�] �&g�Ѫ�Xd���4#c�g��XK�|	���\yd#/B��9����� 2�'Q���v��]���3OT����ޕ��q��Q5�d�Kd{�/ qH0!E��}+�<8���C�� �<�#k4DN��H6�ѱ66c�)}�gP��Z�x��4��Ѫ0)��|g�t9�)T:b��8jN���f	9��:�Q,���+A�v�n���k��R�ɝ{�����e���P`(�RF�P��董$�ѝ��u�z�~�
8���^��@�C�����o~��9��n�����~*{gg�j�%>$��@ �M;�(�!#�NP#��f�������p��k��Z]���N1ÊF�4���X�z�Q�BFe[F"Vb�k���]D+��
��)/��qS5@f�j	���k���I�%�)X�5�����}h��*r|�T&g�R�z�����-'V���F�AWiu[&��d�8+d�y��D�!�~�7�0�������t�.�/�����$�~%Z���$m��"*��U:=?%Y2 S��pl��N�v�O��	Y���A�ŀ�
�9HLS����cmM�g�������#�B���l:q3��d�A�`?G5cg{��qᓏ��w�˭;��U�0 ��K/��4���/�I����|M ��/_���.��hc-���Rm4住>���s��a�� �ʹB�)�l��Fx�Z�2���׻y�&�׏�Q`�Y�9�S�h$�>}�s�X�(����ҽ��ƶ~}��b�r�u����E�b�_�ap�����8�4[o�3��KG�'�qe�Y7 Rӳ����*��AI�K>l��O<EY۫7oi@�U��EVC�Mc'o�B��u�������x�п�ؑ���u��}`<G7�_���mII3��FA���ۂ�����?ן5*R�L�������.�Y/��4�ҿ����!��P�L�������j�9 ���B�T�aԏ�F�H_�;�UC�+�m5bk+KrgtDR1�F={,R�y�d�fۛ1\3���G��F��9Y[�DH,�e�%>��z��]Uö]���c�Ԑ����!�8�dc�Ŭȕu�m�fv:@oWC(�2� ��Yf�"�Й���'�od�l;��%�d0�p�9���B���A�A��z�;D>b͠�a,;�� ��l���6�ѯ��/�O[�Nv(2- �Y�ѡX@P�Ӄ�z�*��˲�]�L� =�#�s��<#$m��4�$-dnn��k��Z��)ǆ��2wĔIc�3z�x��l�3&�椼���p��;��G
�d�&�u������w[��!Ԁv��k���J�@�F��5Z�|�	g3)f鐍E�׃9xO������k����{�h� ��Xf��ֵ+�P�5K?�9*6�?�� ��?�����֛��/�ч��KU�!� �mZ^�N�ח������3G����O˂�6*kYݻ��|����9rD�w��	��pnXA�
'?9=#���o��Ɍ�y�ǕkWO"�Fe �E������?8v�(�ςE.5�H��=�8�Έ�{2���,������A0�֌6��N=	ؒl<	��v�8�ב�99|�(ER>�v���W��9+�AՈ���/�}W������ʎ�KA�{ ���@�̗ٔ�U�%�`4�e$�@y��"���R�o|��kY�^ssYں
YG^z�y2�ԥ.�L�{����o�n��ZC����t�6��ef���3�����`������uD�s�ܬ�̎����2U�K��nD��>#d��ȌV�Y�d�����A!�z��]y�Ïh��`�B�W=&������XY���2?5�6+���,2�(Τ��K��ЂF�w[���w��qkq�Ƌ�0�>/�23��>�����X֑�*���(F���Ѐ�R����RԌT'քK��-�&���l���j�$�@����iA�Z���ZE6�We��V3PքNx�}QSڞ�����G��+t�h�HLjT�絥�������
4�פ�j=�l��N=ϊN���^W�x���20�ѦL�;E�#F��v\���YVO�	����/����*[���L�NA�ĭ����{dsyU3ԊL�ek�˾5��
�C��g����Y���8U�%2 Ǒ��M#bJ�8 O
�!�][���{he �>�ҕ���L�_�)�>zF��{��5t�~��Ԁ��﻾]�_���u�{�L��Kp����� ׎�V�}D ��!�>s挜��z�Ј�X�a}�5y��Sr��q:]���ooo�þ!w����Çd������u�=y�w	�E�O�YY__#�n�P�����D����}*�7NtĮ7OAK���͕e�X]���6�)�J��	�����ɼ:�����n"xۃJ�P�zc�U+V�����u&`�oC%���?1������84+bGt�T�'5*}��L �SG�Wo��7�K6z^�Ҽ:�	�f{j� �qط����6�  j��#ɦ,����F$�����[�r���F�%����G�K�H���k���bF��v]�.���Oʣ'�K9�IZ_<�6����w#*�a�y�h5�jLR�y���@%�`"��Ϯ�ǚU�=����>5h#�*��Ԕ���#f��\�i7X�-�� '���(b�X�v$g��\��Ͽ/��x݌X���@,��qR9��H׎U�B���bc#1E�m�d�߃L���C:���\yL�hB��7��YS3��VWV5���VC��A�i2h�s��ܾqS��j���}
�)~��o���v�ݻ���wߕ��U���;@� �0��f�$U��+;.�(�q��:x8t����95"S-�"�Q㹹�f9og�Vܷ�ny�Z����yxd�D�#�30AP�D��{��`*
i�ְ��� .���L)O~��E4�眎���p?�tEv�9K:C@"� ����X��������;����>�b�0]H��㓍��mnȯ~��v咬�[������.]���nJ���[��4sޮ�o^}C�}�#"��ݠ��E��!C�]�N�9�Ν;��[6n�=�����i�z��T6��������-�	q��Z�t�l�O��W������Z /?"�˚��^Zյc�aPR��+�ۈ:ۓǎɋ�|�A�TQ~G�Ө7eemU�xK��N�`L� d�+t��3����Ou�}���Yz�0����~<-�#�Ɠ>z�埰&혤"`*����~�����жSqI^�*�D�c]��e[޿�7�[B�����8����x��ԼL�SU�8��k�R#��S�U��?p��I	"��	'����r�\ʔRS�3G孈j2�C��=Sey��Y��H�S��U;�����Qۆf�eL9� �fS
��<u����ˉ}<�0��Nr���f�Dփ=jh���*���H}M����<�&��@F�P�5���`I/�����T
���D�3xѯA�Ս���A��s*�����<zr/��#p��ͺff�Ǥ��t��`W?ϒ���7�gѐt�R�b�� ����|�d�A�Ͷ�Eʶ�CG���FO��%�@����ԺܺqM�ݾ+-{�Ō���g��oG�������3\N��ϯ\����\�eS\�����1�Rz_�0�3Ԍ��i��6:��S����Y�q������b�X�^gG0������a�ݲL�Ul{hA�hG�����Fa���w�Ya��zO�ٌg���/�P�âfz9�����}����]V��쬌OMR`��.6��{.�B *r�+H*8$$����ق�`� s��A��!��J˶:����t+�z��?6�}z�>�dDa���^���a��;��Ee�;��S���r��MY^\f��� �zl"���ԁon�����iH����U4�ugIH�C�i�	rY�/9)��R\�*O>~V���濖C{�dcm����Pg<���'N�xiL���Aya<U����(��\w+�weE�}0�a��e(�R��yQHJ�I�(q���"�3n�,��C<M��}�.'&ޱb��!��3�M��E�������ׯ�x�п�v�)�*c>�9��QH}{S5pM��1&��� �.�^�A0h5�w����4�����A���� t�}nnV����XG�QU*�<2�e�����1�mE}��_��|������(P�8-[�ؑ�o�?�b�F
�F����1���`=G�`C�F�.���j_7v��+kr�w����읛~�10�`Lښ�8�!x�b���!�jt,#sS���������\~{񊄚Jg݌���}i����M�pp�*v`�������-��P%<�i�T�N����q�4Sl�=G�\I�e5r���z���zE]3��k�SD�裏�܉�[U'l���fqr����3rg�\�}G�
�7#�(��#��@^yI� �>��<�G\�ɠu/������,Ɉ�ù���#BK	e���>3o�":H�sb�l:3�����Bf�A\.G����qNL�� ���"p�>xH��o�]aE)����4�r� v��,1�hG2g��u���>$���H��o�I1�'�0���~�"xr��#���@��;6�N;���;�cG��p���	鄁ntL Š���h�Sa�M�*Q��#[!�zm��PG2b�����o���E)�����,޺A��Jt�t]=��sr�����˲����=�م9^�������_0�)�+j��>���1��;�7O��n������� 焺
� P��l��K��������8�x��]�?�Cׅ�9�z���8L��� ��~�1�$ KZ���y�/�)���jZ�̫5W������ڲ���V�@48f��j�rP��X�f��M�r��X������3u�����F(�i&���/�T���:�pP���(� �h�3�p%��Q}��C�×�!�Ŝ�qn-���K�ɇ_T��&�zp0`�Bf������c)`]�Z�ܖt�D�Z�jzwF)F6Ձ���������N�s�)��M��Aɉʅ04-k�wdzb\�x���K2=]��G�O�W���,oV��N�e򴗺��%�bc��4��Č��%�6c^|%�Ѝf�$Rf��}[�����C����BV��v_�Æ:�K�0��2��DƬ�g����i��焬r[�K�z>���<%��J���S/7%�7&ծ+-Ԭ4�x
�p@Kez�ۑ�ŷ�\@��nC���=t�j�Ȑ72�+;"9�0�3�o�F� �1+�iVd�(#�[���h�����M��kF`�	����<�O׺#wW6)H0&E8�(�Kýo&�vg� �@��Ɩ��n�`��L3XU�� �8�g��D&<'�����YmI�^�F��iS@��1od�P�^!�6b5��Ν��v�q�'F�l�@y}�L�yu�y6`S,�=�~�s���K�w�:��o �ڕI]??8q�T9̔cd�JL���#nj�t?�M���ŠA~�~2��ɓ`.9���>)�s�}Fv�<�� ����g�� �������A���|�տ��šG++�n�Ӵq_x��F�s���m�u��%��Q��,5uW��~��A5��-�G��R���ц���c��T��Y��f]}��e���E��l�::�F=�f���3��zGzM�B�DybL��A�#�rY>2�&I$2���D8�C����z�Ǚ�^��<v��Wuӌ��e�DQ��ԓrxz�s�fW�;������r��mYZ[#E��nƂAA �t8��22$��v�~A����hv^.��^E�ߣ�ʬЈ���_]Y�ՍMf�@P���EV9_&'���+!0Nb�M�����!��o|�y9v "�'{X�+u���s	{��!<�ic٘�C�5Kv�U� Y��0�B+���!�٤g��4�rhTA�TZ��YmI#�4$jW�����cgKZ�(l��N	Bӽ���!5�@�74	d^; ���w��h04Q)M�3~@�nd���A~V�vNj�-5��e�&�V��i?�t���4���6��p��Y������'��C��kJ�2$�p]p��8��5�i ��=�M�g>�<K�P ����8�&	^H�n�W���^{��a����d(��2�<0"*p�AUD�'���v#4��+
�$��M�	�4��l�9�/�gٜ:�l���&ـ�0����24���`�bBh8-���p�6�Iʔ哹�X�� أ���%�1�D[����>�K����!�|��8���AT�:T%�1�ƄH�X�_�Nr�������R�U�o����1R�5&eu�G�v��DUmw�������v��3iÀ��(�K��0��#�pу4��8�Az�ygV6'[�?�S��>�v�q���Ugus{6����4�釶D�����d��ad���������e�*��N�����墤W�����y�� X�A�& (=8k(�eJ�-J*'!P�VZ��;5�>�3-0�E�]����Pw��F�ي�І�f��`��^�%:/���as����e	��05��4��vV���>&����pî\�&?��Ϙ����v���ETlu\!3�raR�ٔ�@�3�] �3���2�C�<B��<�  �QC���l�����7����:��p� 9ub:��jE���������[���Emu�d�[;�W�ɦ���/�D��S���o޾(�Ŋ��&�+54<�9W8
�B&6�(�	����IdRZ�����<h��q����Ј��9��+��>'�O4��o 4{cl�@1�)@U$0��8��L��']m`��nVD\��'�~x���GF4�9��,�֔�ƭ�w 4{������E`�FIWL Bc,��'�Y�c�<�?���ߴ���:R��P���H'1{��
��[F Y/�-��]P���]oh>e��R<��{蒏M���P1�x
�/�rf'%k�Q���I���	��!�/3A�x�D��d� B�=BF��,d�2�0��h����R>M�����P�l��*�!��s�D)�X�^`�6q_���lmv��r�37�!�8�4�T�K}PAv�j��H!/=,~�&[�+�T�	>���{�5������s��l�"��|scM:#:�D��3	7B��HZ+ɑIo�wK�L2����3��Y]ѕ�i`��$�q�l�VF�>�`p��8�A�f�9�UO����/�+��W���N�kJ�N��(���H�:HK 
�zZ��dˣ���F�z�H\�����F}G���f>�����y;�����wt����H�n�����Tx���p�����:���@�~lOC�6%L��sf��}�DY�~B��͍f��E�
���\�4c$�(XB M�b �,��dj�$�?��� �XY�_�vN��f�p��ۀf�t�2=� E�F��A6���8^�^��^������E�����������0��Kc��'�񳜯�kW/�M0��3��O>c�+�9���f���4�fNI��W�˛�}G�cߗb)'��-�~�E��-5"ٔ-�n0�5�X��ن�*.�s4��]��� ����O��C���3��i��`d��׫>��.��5�I��A�TW(f4c�������k�4{��꺬nnIO���;��_�=��� k�P�um�6}��҅�^<���xsu�p {�r�C�TP��H�j��b�kǹ?���Og�����cNn��ƪnF�ϋ���O���� u8@�/L�i�8�JGFV�gM��3k8 ?Gb%�̱#{���C$��7|�ȶ#;���v�]��������{0cr�q���G�zu0��k(%3crp�>�`A�gfH�J`d�n�V��z�s�5�@Ջg0ގ>�J�Noa�j#h�A��A�ȍo�`aW���=�Y����a���d������T'�nm��� 6�	#�c��8`��K�L�Z�������4:��B�)�j��%�I>'h������-�� ��b����`�0��㸚��qb�������k�����Ho��7�������c��v�j5��:�V�'P
�)]ȑ��S�����_��e��=BIHu�V��+k�\Ne���=1�ne�W�~�o4]�M���{��[�w59t��0����s멑�Q�٨O�F��#VT#qhjRF�MH�9��,G�"�;w���ֶF�"@Q�C�q�M��BH������:��fz�ǆn����b*݃k�����z�323
&+������w�K��b6V��1u֘m%[�fT�>�L��#���rgq����熄�kVԐ�,M�ͺ�����p � @���`6��UǜfvY��i�:�yu�����ǉÇ����D��衒qO߫��ʔ:�+�n�����?x���Ϟ��s������x��g�JFk�u��:��8803����̭Ӫ�`A������@h��\j��cڠ02��ٙ:QW�kU
�<ǜ��dtzZZ��E@�v����� ���G���w�����ҝ�||{K�mkГ�T�̙� b�,|u~�����fK�T��]�Nێ����ìP����~!3�3	�L�̶���F8`Җ��9��"��@9�ОY�������F���<&��D}J�fP�6t��|���c��k��ܜ]����6���J�C�i%��Y`��50�b	 +�xlm���왝���G�=${�g9�v?(��:H�󈎒K��z����B���������v���sU�ܸ.w��t?��AZ�!X@�&dd��{ou��L��_��h8���s��Ӌ$:r8T/�m7y�5]o���nߔ� �{�Y0*lxG�-����R�`�A����݀��R��o�۱��'��ng�̤�T1�^�2BQ����Q������嘠F�.���#�������<�V�E������[7���7�ZER0�햄���1ND^o���TC�r*_�@���2��?D_�X)ӟ�h�
a�2@љ�6'r��D6�;�/��ɵ>�z�U�bk�LW<�Yo��ah�\7�E��Ӭ�](`�������Rqc4�ld��h�l���K�P�z�K�lу��bUcr`�,��L����鵥!#�N�'y��5�t���Z\��:�q=���h�{�jC���p��:��Tµ-��\f_�k:[���N�&��D��S�>���� �y�����GdD�� '�g�����>vXZ������`�2}f�ˁ��K��L
uzn`��8⢎�����<F�,O�9.�:�V �7F��8��=*��:#��9"��<#W�\"��,��g��s�ސ���l7�~�s9{��L̔x��N��c�$[�!b��{��9�{���Gq�88q �Q:�I�iatT&f�J�\�P�k�����[�8��ȑf�_�Kz�(~F��ɞcg�-��F%|�����Z[�Tڤ��h���I75h]���{[rk�/�-=����z��)��m��}�]#�}��}1R.P5��6�x�2�ss�3�] ��-Ѯ�چU�����X��b9$A�;�(!{a�|�~ojvFF��%S s\��� �vN� ���]�ݷ�>j���q�	�#cp�@s��'��p� p��LR�b/�趃�ߍL_<"]+Z-!�y^�G!���ǟ�Ú��_�c^vV�@��O1�= *�6����I�L&��R�J���hQ�f&eaϴ��mʅO���
 ��>�'f.��u�y�~@��*�3B6�}�L`��>B/��ob.��2j?Zm�d�2� ��2���13A��`�%p�K(��c-t��4���o�����#y�C�a�2?�eh1�jO�S�!=�b�לw�Mv�C�~�VJZ���ʎ�͡G�g)Y�:U�u�ݺ�Hg񎤡ݍ�!6� ��F	˶5������Z@IIM�a��7�Vdd�^q1����؀���6_���@@���Z�d�X:���z� �N;����n�e[vӷ(��v"{�Uo/i�_�������)׺���k�b�i!҈���Q�fu���cV�ՑHD4�]�I�����-)��&�Ӭ��ܼ�l-#Y�Jmc��H3#�̱?�_5�7o-zH5���4J�A�҇4eP����9�m��o�R � C�;3-{'ǥ�O�Y���E�{��s5����2������5Lӌ�A����F{J9��T4�K���ӯ�k�8ל
\�Gv �\<��2��0��ܾ�98;���N��\ʴP���z�,��������5ˋuu�L�h�tHO{��*�8 ;:9s�3�3�c԰n�c�c%�%�V���G_�v1�����5;GI��0���|l���m�~C��&�R�l� p����03�i������A����#���0dm� #74�Z��b�1����f�w�ܹ�%�4윴����/���Y9N�*Q>ǀ#�2����nh���X�e`#F��d���Cv8�z��/���v��2L&ef��*W(U�dx�(�5�~W���9y�܃�\��s�v ��@���}��jM�/�޳ٲ�{v:���9��	%����F�0�]v��`O�惿��?�w���8���%QE�	��эF����ܓw������$-��O�`����s���}�����7�X���[n��p�F�ewfwXSʲ�P���x1�XX�<���i���7u��ry��	��3��>��1� �H{,����5�P��HF�'�@׎�I��,-,H�i#_4��L�z��gdE�C�g/^z[n����r 0B��pdmp@�23�Ā9b�
A��>�	��җ�$��wW�N[X�����7�6�
�Q�o}(�oIO�$�`��ooo�_��2��&A��i،s�`P��dN������(�c=���_}�z\��=F�/*lU�t��)Nt�*�hh����Դ�zm�칓�����|��?���e��;7��ϫ|��ꪄ�.�*����Г���BCf��
�C�Ό�����셺V!�A=���F]�´����~/�ȷ�v����O�Sգu�p�x�A'��A%=M�vt�ލ�����+�����mo��Ά���賳G���G��w�C�@�t��ʳ����<X�;Ʃ�f�srtqQV�eJ���ƚ4�aE����}[7��G��������W~(�����l�����J�d��Y��N
�d��g�=`�MWkrxyY���K��ٖ��|S��6X����{A�������I��Lj�]��`~>��t%���������Ĳ��A��Ԍp�k��"� w�g����(S̃�����V[v�z�B:@O>QGѥ�]�h_(˻�#��³�4ȼfIsjhA�[�/Q���,�Mc�.�[��p���U>�}̹�����ȳzK�)���P�|�lF�:ة֌�г��b5���uE�Me���][U�:����tƌ��H��&�p ��u-HWu��d��F�֔��9�֘�W@��f�X�,ycVJ�J�C}&@���#����q�; YQ�oM�A!���|�x��ia4�A��H9N�@:��9���w����e�s�c}�m��0�����s���{�0�	gR ��U+5��$Um���|����9&9����!��󲿷Cn��|��٧/��c��Q�J���zT�ߺIb���u�p|���@��ȞqD玱/��;q�؁�t�8�ٙ���S'u_���͑8L(���,�k0�J�P�RV0=v8�eA� h{S��f��B�i�rJ�#G�K#�����y�_�V�T�(�A�/�C�D%��_c耒�+�{��a'�z�Zd���7�駟�&��u�3�Q��~W"Y�Yh�Ie��1:bo?��`�j��B����F�^���Wt+��a����y�����Q�s�@��mً�`�/t�ڑƮa�M`��~����W��ڏT�o��V��B�E�|�]ȯ�ZY����v�`����8��8t=�Jv��޹���V7�d� ��#{�~�y�:ィ31	6u6 ��Oh��i���������N@�D9Fp���\#���Mf(Y�Fm�gXY���mjG���f
*q�ҟ���%�tU����Y���ȕ^T}'���zE�[�Ծ�y�i�%5�V�1_���Cs�?{���� 3e�,9 �\#��m�~N RwB�"�	HI��|����h\�̌��y�2&�Ha�I����7�ñ�'H��%���%߼�L�JijIV�% ���7ha��8K0����(����N�C,Â��D14�7 �!��lL�\��~]��R[m��膌z9��4Zh2��su��vJ���.4�z��e���-[j֫4�� ������9�A����f&d!��6F6�SH��C�z��˙���g��@����=hC�$*j��v5����5 �Z�U���:�i��:%tG�������ZmF2ך&9���:���{ˌ��z~nd���>����ĩ�������|�p8��q��Բ�Zʧ���z@xg��M3T�y��Y��P=����CB�*�`-���#A�D�ט�_���{�zsg��\ ���N��]���gXk#���AS\�A=��1$��_�G/�=&S����ݻ+|Knݺ%��ȑ��k��n꽶�@�#W����f�|��,j�Z_��9��ŤrϞ~�U�$�(�_�N΁J9�^�W��X�=�mN�RD&4�^��^~�]����̟8q����s�v�;�=���>"����c�C��o,���劔ヤ�U����Ǐ��_�`h���-\ь���;T����*�ыQ��&�k���'�ZR$][��gw�;�k?���h+B���YX�=�[g7�Ԡn�EA�����0H���r�C���R�3Z���F��8؏���uPY#4F�b}�#�aG��{�'E8B��(\!4 �Ue2"Ǿ���&)�"֗�y�wZ��At��Kj�>�h�?ϋ��)R�Y�<�`#Ȳ �(���g���j��
M%�0�|t}'��n�D�i����+�p<�}��҃{w���յCIƛ��4$�:�r\�B���׏�?����p��p��f}g<�>а�G�n��'���(���NBP��nǛQn���eE���{�J�Q=nj�%�Q��j⾤�����BiQ��zA�I*u=�L�Ӟ��`��T�f�A���ؘ�$%��G ���)9u�)Ow�4�׵��9�(_~�9f;@�2���H��6�Iaf\@�$��)q�g�sв��n�m}v�"�'8��f�(5�ԧ�!��"pԥ���$���'�����(��w�%s�^%�1�(055�bgu'jdg%�����?G�d�`��B�A����2"�}���f���sfX�V)�}�VG�v�t�$EqH>��H���fۑ��$�>�l�l�����:ӎ	�`6z�S���`�@\�7v�zz�
L1M���
�s��6D��h�1�(��3�M��}�P��Me6��b���*%�]�L\f�,H�cаFq�k�����q����X[L��%������c���ʐ +��679�pїh�pk`�;���E�p�I�
`6�d���妨M�Hg����ލ�7_|�9�6�i������n^���{�\�XC(#˄���*���(7�U#�q��[��nӰ�'M������ە�g�X��:��i2��]���ޑ����2�ptp�a��KYކ���'<�J��}Vy����_��T�{��%��O"��~�%��9_>;ұ�a��~������쉮heܵ e_���`���jb���
�[�`N<��9�Om���c0\�5���PN��eP5Ijc0�����A	.���sKe "�{�^�vDA6�ܺtiQM�%G��G�*/B�%��ߙ�@T��y��$��"N*<8a_�*��;P�&����H�:JոE�@�q���߶o���s�O��/y<���`��ݛw�쫡�iVZ�j�c_��=L�%X�Л���V����)!�G�#��,��(�"(@��h�N %8唭 Z�*�V�~�?��S�U�՛z�wRʚ��>tA�!W�`8ir�N�G,��Z�g�R��O�����f���3�Q�2b] @�:�C�B�k���(	�a#� �4�?b����Tv�7I��ȵ�� ��{��+���s�[`Q��dWǎ�Q�Kˀ3R��}f�@�B�N�.����5�[e,{g��4���m�i�D�Rq���`����t�9<���W�C�6s�`!p��*��0V6�l���G y�h������Y8�,��]ɫ���9�<�w�e��IY:tT6�7ܸO^�6ÉYa�c1�8cn�{m�*A1�f�=��e(.�Í�4@i`3θ���I�"@��$j�����=)-�0o�5 �Y�G0����ي���u���VH.��5��ٓB�s��˶^��b��~���{؟*@ � ��ؼ$W�Iw��}Y�s�]��� ��d&����>P�[���?�chٜ���(5��>4��:��� �(�l�G[���L��f�*T $�-��:�'�PE/gYڂMa�4�BǇ>uN��&������K_}Qi���3�o˭������Ʌ���9�|�h&ϑ,��LVW�-�f���?��)2��6)���ޑw�ݤX��Ɩ�?w��o=�3���������Hg�Z?��U��Z�*�_�6B�3 Y��T@�����*/��E������#���f�u�d� ����t�	�(]��iغ�8G�s>��|�����L^�w�jl�-OTL�a��8�ƴ;b��L���\�y6&�A)&n�����ۜc�O�U��A��a`�A0��ո|��m.����� �1𒟝D���
wn��c��Ώ��Q?bB
Ǎ��Ŝk~�p��:�
�z�=ҵ������T�}��K��C��]���`0S'�Ԍ4u17 �P�Wk5%hZ��F60�<|��iJ�r�hc�0�F�LiQytV��� ���{/.,��5=;c$,Eq�Z�����N>���ݭ�����A{t����o�m��O�{��/V5����BU��Y�Z�ÂJQ��H{����F����������v$TG��ۢ@��yi�>�p��:���sY�wJz��2�F���0:���m���`��L"�sB���26 ��Pm�1���,��3�2>$�6�SK"cj��	��"\'Ɛ���6+�����͎��dmu@iJ8sP�n�l���
I<�i����ôZ��}$T��s&W4���z@�;1�`�5+ޤq(ܿ�q������8 ]n2p����U ��t�6;����7��#��+�9���3�{>tL��������BU��Y��鿻[��g��u��/16���F|O�zCW��ha!�笜��1*A�ް<��vr�>ȡQ,	Y}���i]�
dk5hAv��k�"��zn�%l9(���N�<7:]~��`ǰ�!�a����~W65 �s�>(p����3��k�����,��E�!١u����gO�K_yQ�f8��W���;���,��M�D�������2u�P���  �y�~��!�Ǵ�k��ʌ�)vΝ;��Ӑ��>��Ğ�~�.i���������~�>t�
�\L���7[�<uR��,���M����K�jE�ӐDE�}�5���u�Ux������uy5B�B�lI���N㊵)q�����a5��l���L{���2�_��*���&b,yC��}��"�����X{�6+4f���'(�L��kd��~ًgG���re�f��[!�Y:�qe r�a�2��?��u��0幕|	NC!v<�$�b�3���
Y�B�Z��&����0=���V�Ň��82��2;;�|�t��th~^j������b����Y�!FO� L����㠎���0S�RIF���`=%V��^A�ȱc\�� ��k ���C�97�湶����//����]���B\mh�|V�����o�f��,F�t�/�H�eJ�}0�5b����C���%L�n[��� �k}�4��d׸f��5L��iW�MG˱��4��@G���5�aSҚ��Y�$������2'*�@)8wdDI�2M1��)uđs�9���*�pL���6>�4(��ݑ�~&{z�[�1�YH�����@1jjZf4 z��m�j�,��PY � p�����qe�Ǡ���.-Y��c[ޏ��rC�R���1����3�ܯ��
i�u��I]�1q
�xAd"d����5r�< �q2��3�\{"t���ͤ�N���g�O�q*8�Ԣ~�"Y�b��vQL<�F�+Ȱ&(��`�Jg߰ފǙx�SR�z��_�ٿ�=u��؏�qK��C@�2y�l���$�Y��,׷-\�c�5��$�� TK����db�eg�f�<EslR�b�|��ș��48���֦\�zE���rT�u����k�����c�I�N��FÄNP��yG��<����k���@�5:��&$L�dSC[a��@A���5}��D�!���]�y=zX��XQC�I��Nq��5�_۔D���׮Kx㦘���H�������|��f��6���S�z�x^����T�Ec��5؁}�1mNG����7bP!Aϙ�)�¾~΂�p��̰d3̛�����б��UÉ�
J�G�O��`��ֆ{擸�q��r��r��/eL�b��2���������m�~ȳ|�n����e�9�����ǳ�+�T��hbc{G��ėB�Y"�s�!*/,�`�����>��ǵ��A;�(:r=,��C��I���h�׾����j/ݻ�ݖ�T$��eW���d��\�ey�%
;�����,:�mfu��M��:r\j�D�e�Y�vw����Q>����nY�^�YZ��*�e�X<#:Qd(�n*���x �liB����g����Mi��Y䭟��S����{�C�I+6/����Ȃ"�s'va����P`�+\9\�aTc�,��(��Z<7}�N[����(@S�l��,��b-�:(/Q��ە3������	��OP��=�\*��{2K�ܜ��|aB��F���@�?bo��iB�4M-[��5�ː�1@���ў! �X��?+��6~��-�j�G�H�K �?ÔU��s�j��5�f��]f�6Rd$�3�7�U>c �"2�Y)ְ��{fm�8��G���$^�gr�0� ����٢�1�~zAV�5��[w�Ӂq�9ֶ��c�n��M��c��KC9�̌Ρ�sw�,�Binc��z��r�"�B�I|���i����W_���>q\�>������ۗޤ�+Z�D�Op�{�����2��R�>5��z3$��x�,}?_�B��K_�Gr�������4Ѐ3�����vMb-�<e[���S�N���4�W�/_���oɉ�%��]�����	LO��|7�;r��-sS-������Ox�]�%�ֿ���</A��F������,�.]b`�s�9��F����5�w��l<�+�n�zl�麏1���#�xEB#����ᰒ�o�L�ߊX����V����dF8Oi��Ag�r4�q��=ȹi���L��Ɂn"�հ����'�u�%�.�B�|�QrHޑ�� ��C�c�jM4��0����},�(E��t�8']�`�`˝(�07FO;�r_:��O�����I���$�+��cp�#�u�Ӈ��p�7�SH�)p`��S���(�֩��R��7#DV'3`��z�@k� ͒����uF���V茾�nt��,q�B���A1�O�@�ǖf�MͶ{Ֆ��~(��D��:�Xo��C+DtV㌠�k~(�o]'X�ޜq��t����f#����,�
p�xH(�1���֐�V
A� 2�3�s�#����s������W�{�}f���������$ڀsG6��G���� ��sg�0��ӌYCO�s3M���z��\F���d��h:퐭�<l��������Tǟ�=	�����cF,��?����d��B5�;j��
ZD�s�ݬm�IP��_#ʁ(��h\0r(|f�9�q<f!\Ϲ���?E����W��O����3Y��#�O˦뻻7R�-�0��0���;�q�W53d&h�d��y��*��u�� `����V�C���%M����:;:a���ڭZX�e��� �j�ک�Vv��AVf�>G�T;��_8$��(t*Z�e�x��U����2����!��A�! �v�J���L������&�^=-5J�U�T�kM9���=s��;0������~�Ր��e�x�qU3ȹ�L�,<v�
�o��s�d�?�[F�k�nYl�1�@��Q�������.�)ͤ���̨�}�K_$�Rgu��+�ё������^�^C��ڕ��z�I�j6���db|�5[�ʕk7�h�X	�� 1r����U0Hm��Vi�˛����g�&�N��1:������h��z/D�Հ��İ�O{P��W���~Wu_�R����@B�1=�GW�����������(*:A0�b�L�[���� V�a��O�Y��v��fFye�r'sI ��=�i�Ja�UӨ�����(*AV��VM��F)	��W�F�Iutq��:�F@nV��ԛ�(m�s�>��? �
�Bm�B�xn(~f�O�zo��u]'���u�н��.A��(t3��٣�z��A���{�����|�3�4 ��(����1u��@�fe�^u"e�D8[*�B�������;d)Vn�r
���s�&O�r�����"k�6\+�?�C��J��d�ϤD�SIG�pG�|����E�]Y��ԙ�2��捫�\Q9�ZUG^�f�4�t�ƈ@u�f1���H�Ap����<g����AN�b@��c][]%��S'H���Y�����{�[�q���o\�)۳34P@�~|�cn�9 Џ�q ��t��X��h���Z�B�>c�?�!��slgu���+�Ge�3�X�g�rx�c.���U�P�L�g�H��R@�M��s���\8w^jCֶ��G?�� � e�h)�6�qY�F��w�׍?�q���47���-�>�x,+J��f�� ���ٗ��>�!�����̌R�һ�É����t�pA� a�>�:��j��<���f��z_��Ʈ��7J���
J��q�����ht��d���i`�1�WJ�jH�1��YJ�"�R/��"�=O���tg�6r���P�+������!U�R�������gu���x�w�����C/|���P�Ԁ�x�ݷ9�`�Ԇfo6�%��;/ުȃ���V��?ޕT'[:�\i1�E;��a4��wok�~���3���>y���;�!��I4�2 ��s�^w~(�>������<{���j�t�������T���ٕ���iu���;�c�>dl�Y�"b�����"%O>��D��,����U���0���}�ߦ �?Z���Y�`K�R���Uvu�	�-�8�'��׋��������X�#��ڂ�O�W|�[��'���q#�?�c���x���/����������E[�f��$��	4"	0G� %��u���z��Տ>|�|B��á�ZIv ^X�wD�ҏ�����L�s��m�	%l���P�1��� K���������?xd��0�c�� �[��V2�!j�7���?��4Ԑ�<�o\dyyog��V�^������D*ͺ�-�LxVZS�כ��3�	;���Ao4*H*.gdِ�� }�&5"������=y��7���#2ۊ���3��o~S�]�JjN�s�5�g��YZ�c�A�O}���Mf��V��x�����Ц�K�Ws�X��`��i�;�s����Z6���5fT&�׹�fUǗ4�ɥ6ؕ��i>ۅ�i����NI8�� YlM�7��os������>ؐ�7?�a�e��D����HfWv�k%s�+�dm�������d���{qNxhY�K��l;$	O6�̒*����D�"R�VFK@�$+㜍4���2Ώ}K`П��\����QjΥp�cT�g�����	�����N&�x�������O��K�@O���M�Qw���I��k~ϗ��k�=�.�X,<R�z��3^7F�p�'��`O=$'����7�Yn~x��9���Qb�������)�z����ۨ�&erj�{�k+N�u��c��5�`�m,�I?pn5��O��wtn��s��m+�0R ȧ\�{�[	���>��g�ܹ��ݿ�����op
��o�[�'g.<�??'�޽"�4�g���J��2�� Ј6ҥ��^LT���-��Y�$�q8�sA�9�4�"����}B"��������1ɐ�Q��`T�4��?�����y�'�_Ώ~���'!�8:�KWo�H��̝S��Z�C'Z�(��k��*e��cɜI�G18�����d��� W�1���GT�Q�sAX���s:
i��S���&���4�T�R��n,/�3�z�?*zFz]7�a�R��<�VQF�bT
0(�j��r����YJeBu.p�hP���N�����a��K�}FV�}B�fU���/ȗ��e��+/3��&��Jλ�]��{��e׺?��l�����<����e__���h\}���+�r���A�M�_W���&�"���5!�X0��I�:��t�4#�k��̼4�g�Qf���M �H��W�����3O��X����`�
��R��L��(;O{�V���Z�I��Ɨ�c��*T�F��=�=7i�Q�9����B(m����Ι��֢����/��#�'h�W��Ni����z�`>����P��:{���{��qLy�G�Jyބ�p�� %�̏�w��6@N�3�$"b�<�@:��u���P5����Q4'n�ܐ���!#���6��<�N�j��="�91�?j���:<�Ad���mr��Ȟ���&Kʑ�L=�>����Hꉭ@8��z�>P�i ��03=�*�.fށa&�;"Ο���1 ���K%Ǻ��<ӵ�;�K���r����}�j�J�o�����˯��ֶ��pޑhY&�6&���14���J��t���=��^�q��tL�����x//�
�r���P/�F��	�͒5�OT��y�t������B�ǧ�/w<�.:�i�JT!�I[[���_�)E��y��F��q4Q�+d���9-;t1�9�BDڏ���A?��4�0��廙�,c��	hߞ:��l�X:��lh�VM��ڔtv�5�d��!9}�̬���|�Ѫ������+@����!ٺ�,�U�@2ɋ:h��C�;!�&������>uB��1����{����������W��ex��a(��$a�0��^K5�I�ըX��۶���������B��{j��#7n�IRk�T%����?�uS�V����{��sSri�-����=t�4���<���o��q�k`s��-y��׬h$�EC�z�U90(96Ofc�>���A�U�Y1�,�~���eR#A��Y8h"ą�p<�z#���Q��-BVR@@S��kȉ8�a��
��5md���L�of��<G� �A��(O��'��n����Z��a.#�Yr�����"g�c
��y��g�s����V��x=v����K`�{�����5't6�����
�F%��E9s���L(��pn���׎�r��66q���7��8E��{�_as���94/�{��և��N��0�:�V_��%3��N�:'�s������&�td<��@09�4u�x���No�@C\���;����U�?���Vl��0N�%>�A��F��g�a��� `2���u���}$�#0L4�A�2��BO�Q�&΃����ج$�(M��t��$Z����D���8��Gw����	 2-cj#��u�9��)�B1� �zo�8��Łh�ئ�:r�G��a�Ǩ!�h����Q�L#td�7ʰ��!U�*���� -��k�0��h5�饺:vJfW��v��Y��_�(okv^�(���U�C������͏"�a,
s֚9�,��eMo����;ߑ�VS��7�.5�@�.\�?��?f��7ߐ����$��;��`/5����]5t�qK�k�8���<��~|jwХ���	H{��T`��npT�-�����g��N=.�;�R�}��fLUY�]�c��y}�s_��_���9�΍��������af�p��q=?�<;��N�g`02�1�%�t��Y32b��>��3
������A�V	HP�o�c�sS�rԦ w�t����c�Q����h��׆�I���"�x�b��~�a����~�ꀸvA�WU��L.��S\_T�2���S�+�Kĵ21�3��>i�>=�&0���s�n/�]�� ��u7�M��3Osk�w�}��� 1
�d�!��f�r;���bP�	�SsU��,v)J������D��v�UG���M�ԏ��(Fږ�����5��ρe@Ђ@y���٨����)O�:����˗Y���?$_�����|��Fn�-��Ɖ�|T�� �G���5&2W(�ܾ�>�{���g����u>hb�E�{gPl#k����kVa����������Ď�'�B��mV�_�Kxe�m|ܘeV��K�ސ�2F�
���s�41J%/4A������D��<�z��oL5@�H�F� ��ƴf�����TkV�:6e�ʙ�%�F�d7�e�������Y}M"��;�������{r��}�QcUiV��Q��fM����#3j�|0����k4��"�ń�2Wȷ���r��qy��Y�v��_}I.�c���J�]y_��� ���N�M�a���r��k	��PW���(� �g���DT_9���Y\�!M	�t*�i��M���b������}�i��k��ưW�_~^>����Y��^��7���|W^��kj�)e���#xh�Z�0J�8O��e�v�HQ8�`��ǁ���T�j�]�'�0�*�X=���:O��X#�5:��e�s���T�Vf�6Ah� Nժu�f��
�r�cn�]����&��/(���$'�@9�o��1
C���8<�;	���>�7~�w�lVLxnG��#��.�G��	��M�Xᾳ����;T+��124:N0�y'TC��^+�Ľ#�Y�8���ck�M�;?#�b&ޡ{�+E��mu�ݵ�f��ѦѤ������9�&���=�Թ������� ��x����G�Yu?}萼�A��=G�z �0��Rm��G��α8_YvMׂ����P���%���Ev����.�hx߲����:AU�8ab�9��2�~�'�:C�(�雘�e�
d�?=>���9�qJ�p.ʟ ��F\�N���1�Mm,����E�ހ�E�R%�=CG��z0�36բ�|���TW�(�C��k`��D�-2���~[z�>�vZ��l��}_�85-��#'ɺ���ѧ���f����v{_�4�F�wv��	10��y�4Xt�H�����Gϧ��w������_���/��ET�dvnA~���=�ݍ-"�˺�"�$[�~4��Ч��r��+,��������R����q]�E�B^�կ��#�l�Z2 �
��3=3'��2�?~T�}�554�4j-�!k ��'��ݗ ���J^}��,��I,[��*f��j�,��0=p:Z�9��������x��x�Nv���%q
�i��[S����2KCV:�n�Q��zq�T	���� B��p��'}k^Rؒ`8u\GVV�ƇW(U��t�Ҟ��•V�fe"�+*�#��:#�܂���Cs'��x���('T
��8��@�����~�7_�?�BGE+EYe�B9�0(��"���E�*����al=4A �Y8�v�FQG0��d�F�o���9ZؐH�%�I���2r�����E�)CCK(�;�:���z���y]�΍��$%fE|��{jjrA�,f�{��8'��굛�}����ɣG���h��}���#��W�΃'1nW��ڀ���v� e�c,�پ��:��y΀��[���d��{����<����r$�F3N�$���X�G�Zyd���q�x,(w�����:ّ�������MF�Grp�����(�و�#b�#����9������٣(	<���̴nژ	� 0۱���Ew�fQ���lt�)$�r}���R�C�@�5ͯ)�R�iJF�1q!P�Я�8[��TC)���q�kbN7�������B����o�;���U>����jrb�&ёc�rh���<t>G�`��C8��^WsqY^~�-bz����=0^�!��tH^��oRd���b�Z � � &40�>~��4����%i���+�J��dc����ٿ�s��^a�������9N �D����{�i�G{���P�LGD��ȲF�-�� �s�$���9J��y3�S����AD"�Ξ�qt��{������3zM�N��Q���H-�Y&�}��U)b���"�FV��cZ��k~Z��)ه,��z�)��>�Q�$d;�k�[a���8B�ٶ�F����I�zs� r��<�k��F�<:����3�D��98�����(<�C�4��Xܤ�ˑe�^rp�C=��VEX`�j��z>�Ժ��(�"�לN|_��k�ޕ��l\ ��~����5�̸�c/��4H>�4�鲱_�X`8~����ST�2	��<`�c����a`�su}�v�^q$XS��]��3H��x8"ix,m�k�^���6�.��}r�˂Qư*I#���>ϘR��1j�lT����,�o���|1bJ�sـ��Q�N�l&�r�Q�%瀯V5�������̹��άmn����N�xhg$J� a��l�?����'C�	��3���0yhЏK0Z�}�3(��1UV'����@��v:�X�1	ô����]J�����?�B{�*a�& ���}R��W���\�wbr>4GӃ@T/}k��Эu0`�5��3�Gy�N!�Fy�N�����Ԉ�����?~U�W���|�������n�2�M���0��ۨ4p�:�#��x�)��'oaNO�:7�Q��9t��l�C���ο� ���{sڤ���Óo���4� ��{��w����\}�C��B���7��廙k�>64���F�mM�sT��_����]0(�����b��\���g⇪�ݝ��&����29s��LO5dgk�e@���
���Z��+���qr�<���I�bq���݂�Eh�)�'8�a0���w{ӹG;dK$"��Af�x�Ldx�zj<w2�~�����_R���</��張�R3n0k8[���E��F*` ����&Kב+��@ c�mۯ��I.�3�b���ʱ�363�yb���Xr���lN�J�Y�w[���C�|Ey	�sU�	T�Gy��)�u�IYQ"�Tp�r �g��F����ӨUda<ިBB
f<g�P�N"�P��]:��W/xo���e��U�>�q �j�����O�-��X���A�W�,����l_i����YK�5ˇ�Ȭ-m�{=]��3{���r[�&��N�#ᧀ��p<����\������]$�'�Z�<�����w�Ȋ� �z���G����V5S�}��ٿnF�M�#�|�0�iV��auK�n�+�ņ��2�3wc"׈�D�ѭ3E���`�p�Y[8��i�l}�|�Q6�w�m��^��ܺyE�x�'��ٳ2Ӭ1p �.+
7h���N�$��E�}��vG.����H=��z���U�5������k�&A�e�e�O!�Lq������qŲ*��ekm]�޾#��u�O?.��i�B�T�^�ݖǭ���ڂdN �D)ˣ[�q+���9�"��=���s<�՗,5�95��K�r���l��˽�7t}�m�+6�U�	���egw�8��4�]׸t��\i�g��}�k�q����G��$T ر�3��c�F��8�A�"���O,�B��6"}�o��YX��b`#f�y��������es�B�4���#7��cm�y� ���=��pvo�L�����3�t�%��a%�x�/�u�y�I��m|`1����� \_y�Q��2=���	ܻ��mf�B�r���<7|d�k
�	�(*����ѿȾ�@/s�5��pZ&4�*G8��6��Ɇl�p��T��{�G_�_W}A����L5��RB1���ٿ�63�ֹ�|Zr�������^@��B��Һ12�{�>:-���_���#}m��n�G�3,�<� :�]�W����d�ŲnLG̅�����;*[�Z����� ]D��1d���5� �a1b���i]C� U �0�������KvI{p�gzcגJ>긼g&i(t�d�J���ʮ:��֤c��5�GJ-v��Չ�o��@#w�hw�ž[൶C:Ɏ����R�
�-(��|�@ˋ-�������f�w$�[��S��G��E���;T��ސ��0C�O{=����B]|X,�|�U�� 
����]����ݻ���)�E��%��5:.G�$.k4u��e��e�Pq&�	J� ���[P�v�6����Lsk�༼$>�C�5�h�Q�	�h��~X}��7�Ӷ*�{W��
�������'��M��ysW4����#p 3��@\U�N��1�UCp8����{t�Yq�:~�����^<\U��4x��pf�Ϡ�K�T�ܾ/�]���|]�љO��= ����M��m=�`,��ɧw�G��>x��z$�J��>C\�'cB&?����6W��{�ݫ�����@u�D���
�$pT�e_^?��6�����ˡ������YӠ���Vq���a`(d*�����Sh�?����'�H��a����7��g'�sunv���(ɜ��)��e�7�@gށMiH=^Rt 
�ˍ범0vѿ���A�Ȫ�cL-a�DzoR��Zj�>��Sr����ǫ'U���F+���'�9L��b<��~���qA�~��{��{�3���pY��Q ������Y^�&t�9*c�f�&G[Kr���~��ڦz�P�����1(Ib��;��K�W?~Y��T{#y���r���`��z�q������l	 !��4�By#��0� K��
�Pڮ�}p��U��@ՙ|p�Y� J��V���\-l����Q�h�蓈��=H��_��\o�6���B}�r��Ǭ����y"n��pٯQK�"�!�S��-G["��!9��>�n�z��t~�S�2x��'p	���}��s�)6�g�r��/��k�
�l]	?5�[�e��9� 19�1-2Eƕ� Ka�Ө\-��\Xl�%����\L�S�@�,?�v��D��2`�	Ԭ�L�ρ �Ӂ�7��E��bwf�M�z����E�r�LT�|���F���1I�.�;�)��ad����}��(�p<A;9�6�y�y ����(�f5���e8&*����C�k쑍����á�P�������}YǤ�4xLn�_���z>|�q�,ʲ�����|��^���yX2h9Dl�4%�0�2��0��Q,G{���M9r���Qn� �
��>�ycC7c~8/����:�_{�E�ڋ�SV��)��&Fm��X��:���	��.�^�>�o�8�����Sg��ں<���sL DI���J-����!����C�mE,'BB�]����)�� �!�[�:����h1�j��_���!�X5��+Z��
��1�~{jҭ!hU��Uw���$��,�pMtSe���m��"�� �Q����3��F']ٞjt���N�����8��|/�܁E���k_.h�X��	J(a�S�iƄ���Ӱ�17�@d� ����G=� �vM�4�7[u�:��eҩ��h�<8B���;��1	A���~�e�c�&����É*��>����O�i��Q�!��jb�a/�3�7&�j�'�h���������C�G��}zXS<p�깫zd�,f2��� d8*��X�qe��p��̍:����a=B�D���@Χ�LkS� �Y�/~�!?��zn�jXm�I�u���Ȣ�ևQ�>p���ݩ�G���[������u�U��H��|z|���r��/J��Gu�_�I$1��NK�'Տ��s�����15d�Ÿ�M��I��ڒ������BQ�a�x+�%�����BK�'�#T������;��'�\�+�N���~Ag�E�\(D�ƙ�\$�2�� ��U�{bqAf��n!K�@��T��!�sM��Z��}�ey��:�ew�E�h=26(���a\�'�|� �]U�^w ��u��lo��c�H�d(.Av�GH/���'��(s�]B4|F*Ҕ�k`�����k��~P%���ΎLU��v$W|�/U�0��e1�����@�'�53
2NT(|F�u�U�BV!��t���:��Hh�\q�M�[�9���{H=X��Y�2��
�Ϭ�b����2*�c}r��;�~jF8�X����%�Hv:[�
.�.  ��IDATX]p�p\T4�O8>�g7�:T��HQ[����C�B���_�BC�O�8~�g�
)�n��"^k:p��w�zw��G0��|}�e�|z��y��V8圲Y
$��,u�(�BR���>!�p�B�QƇK�lq���;��L�a�w�����<�H9�FB�އj!\3���^Ϝ=�4SfUn��������"f��$Ǉ!H���8��Jn2�@���	��\�+WĂ�,�x�>y���>8��A0f����]Y[�(�xv�%U���b6�BZTol�����H��Y:-	ܘ��5[R"xʜ�Ѩ�'��b܇�e�b,P��U��9f�iUkqV�֋��FQ�Q�ђZ�)U����H�`,�3Q�~�H&��]�#<(�Ӷ�uq�����@��bFMg�9]��@��n�~�L��=%�ܪ>Z�<,7�S C'6���"�8#��W��A�\|ňX��s{�-����F��~�@ϣ�Yĝ�	��L�����r��Y9v��3?W�\K >��1-0 ����qp�&PB=攜?J���?����˟��w������u��t�ץ��	KԹ MP_�p�(je�p����.�p �<��'�"�I�"S"苡��Z���:�!2��3��2dh�o�yr�`вq��g�f{���NW�������n�+$r�u����C5�`��6G�c5�x�,�B�NY,�pQ�\2�J����'����5�\��(e�'��U��Ul���g�B�x��R6�,숑)b0�r2{��@a 8ҞB�͓���00^��$�@o�뚙�s���we�Q�Z2Aǰp$`ӳ�Ȝ���9۟K6�'�Ӳb��cRz��C����{3�QI`{��bϪbUu�QU���	�V@*���0;��G��QdYy�[ev��k�^7x��
�����w��p�_� ����ܑɳ����X<�w���Ǹ���>8_LtP��U�yF�`�Ba��ʀ�&�*�t��������}��,�Uq`�������(Xl�	��1�̌�k�;T�qc��%:���aD	�v0��&Y�f����iŵ �S]�9Njq�ht8�ُ�s�>q��T`<��k�>�-�O�f>�,���D�h`y)7mL�7��,_ifج�d�������{�� �
�8�PB��Wg	�#��tv�I�ݻ+�����P�ˆ��_oT�6���#j���:���w����89���y�&̷�W���3��wU3�W^yE^��Od��UdqeY6�v�13E@��~�=��M5F�ƃ#]d��tGD��}�K����&�s-�4hh6���qY�sCP�����L#@���Z&b>��F�klVAX�|a��w���=�&�'��5�R�{�<d�`Y? Ш0%0�:� "ɭ
c(a��7�4�TP�����'�C䣒	G�D1ǧ�� *o�R6�t�B%4�6(�
#�+^�&e�9��F��fQ9&"2"���5)�	��<G�XIf����,�k���B��I65�h;����:`fY��Q���4�_����P���r:θ�8�1�m�`�/;TV5����j���M�s�i����4� !@޿Zݑ̌�qq�$4�/Sj�^V���8�)��D���tt�+5k� �hI�b���ސ�ԝ�]�d��S�?|$��=��,b��1Ք���Y�j5����v{gO>�w�cat��������g�}�I��o�-.�9�Fײ���LY�t�<'��zL����3S���̖%zs���CZ�YmO�ޢ��P��L�s���;t����;����&h�=��،y&A8����-+�U�0�^C��ޟ����ְ~�]�����O�M��d?$(�%cuu8 �0]�0jA4��FG3f�`Ik�3A����j��`����ɑ�+]�Ȇh� z�0�}�cR+�?������ל�CN]�n�`�exoMT�e)q���z�PD�5Z�IC"�[B�R�p�4 :�s�z�m��@b��h��4d_#��5%{�[�T#������.W�<���e
�LMV�`(a��i����y&u��1��^���醼��s��0#k��jPs[6ܧ� J���f����l`�Xf"4+$�4��.hW{#5���K
�<�|�9�T�`6i��s�SHǒ�-#B����Ha5e[���8��������2�[0���b$�\@�l2p�֫]���w0�ZK��ȁ��r��ӥ�72Ǚ�9h�/=*Alq��	�b�l�o9��,=�I� ���9�#�_�����2St�d$�Q�������p쩣þ�v��������3g�{���g��4s������@_ہ�.�c��r�u�q�tM%.0���a��54L�{�e��U'p��V]F2� �B�gZ��������Ml�D�Q׀Aϕ���K��ǯ�I\	�~�Lzv���&!Ln�d���3����I&8_�Hz��]�Y=��D�
O��Z�kiTc�K�ò%�us
g�T�O�'|<��rR?[r���I\}m��#&Х��8&��|Y�ڜ�o�ܜ�3����b���Q�YA�I(P�p���Β%5D�h���NzZ��҂,���;0"�v�����Ո*$p���l\@�cͨ��Df�P7ALc��c���G��=F���J�T�|�F��wϞ5��:Qn|P�����C��C�w��DT$RA�N�"����&�ܗ��9뫩����.�!�|}�^h4��c�B��w���'�߃�kj֏ި8r�,3���!"�~[��{ي�������'��?�$ݘ�LxQ�֏R����.h�"�l�`%-���QS�{�6GM3�^�����#���Xh��{�l��t^�j<���ƶ��v������N�7닊�Ϣ���}oܸ!���!+'�թ/�$�8���1E�j�����<M����#��9w��EJ��?!�M���ن��-���p�y8r����t���,�����61&9�ť�$�8"����ԱU�\!Hr���<����ruS�Ë�r��Q7
f�\-�;'W&3	WWky�ph�S�Mڐ�����I<e��n4.�����a��{`y��ڇ[�w��g@2�W�s������`-t����������9y��K������N��'��ӧOS+�7ߔ��}�ƭ6�5$8��7vB?.��cj����e�P�~��S �#9Ϩ,���	ɂ@~T	2"���3����O��������1����"��e��QH	`3���ݹ��CK[d��D�r�(���eƏ8��2�ǈ�8�����=�8�����Ӡ/��F"�`���:�S�P�3r��Q9�?_�L{N�:ʘ�aDD��֭;��������F�=i����p��U
:�)�����Ȳ3�$��0JÅ���A���w�lb8�u�G�eƍt�l�z�)y�+̌[-����4Q1��f$��|�on�J��I�s0�ᚡ^;2+j�gf���mʌ��c�e��/�nߗ�n�]ͤ�5����:wu���RP'�S:&A�`X�ti��|�6x���^g���mo��˗�>)=��5 �z�Ӡ�{��{��IU�C,�`�V�Շ�ߧ� H5�T l�������.���������p+M�	����7��7���n��ep5�]1]��l[����@� ��Fmu�T��$�E� s��pXM?��Ѻ[Y�ęT5���8���͏>�3�CvY���&��>"�K�������]l����6��`f�GP̋�яld�Z�/���G����PE�1eq��Qr��/.ɡC����=T�/Y�GU!v=pW����յ�����|杘wd)�Y��I���<�}�%o��@�;���{;]Y��"Hp���ȥ���\E��ܛ'��cG˫/�,�ǿ�t����yY�o��o�7����ɓ'姯�v.�&` )���Ą_��h��{�_����������&V�?�I�5_1 h�p#{XC�޺$ih�ydJ�O����Cϳt��.���PA0ч*��^:t�ԹO��f���m���l�Y�QH�g5-�-��8͊i]ݏ�x�z��Fv8Id�~����t�-5F'4{:sxE>��Yu�ꜙ��k�Y�h]Q�xd����o�#o\z��.rr�f'�g�����B�%��>�L�8T��R���	��Đ�ab���H�33dwB�}���e�5[rW����:r��7���n�S�j �������������m3[D6����	Y<�߇��P�;/{Ìd4�k���yR�����A���ܺ��l޻-�jKV�DG^~<��:a42�[tA	G�w�������[��/��_�O���f�{R�ƙ.y�D �$'��$U��"�}I*���H�tkJzz�ȀM�$��!ӧ̪^;P��\�C��7��$aOƲ3���5Z
�����΂�/]�`_���W�fx�[����C�,���X|)F�v����Q��VJ�]��5�<?Wbg��b}{8V"��*p����}��r7��MO�ƁUV�PVo���j0���LL���
6Ad�Î��9�P��N����<!k�|P�BW@ꆐ/c̓��CC�|hT���[^/��{��1�6#���?2y+(�{,���3h`m�κ��ǲ��mR�n�bF�F�z����� �l����!����h��̔loo�Zh𞼩Y����os�B@���}Sd�����f�W�mOΞO��=��1��� ɿ�G5��&�D�����wN���i�GŐ�������p���8���c����u���r�G���z蘱D\V�Qs�+=٧��f���CIh�U)P���F�ˌ�pA�|���^I���IQ�i�a=MK҆�6�!�1��%�sǏ��e����>f�y��c��֬ѡ�=vD��H:�Lo||�J����h��u`�B���J��(%����P�p8�
	uܝ�~�:2����ƭ�Q���g>+/|�y#���_\>$UݘW��@�����!O�9a�M?�Ƈ�Y"KP
�� +\��5CQ��t� 8�˳S�<sF�������������)�[�pĔllnˋ/�(�;�$7�:)��U9�rB��[ߒ˗�[/.4�w���Co��}d�Q�lvT٪�����}6��i�����75EH��s�V��z���bF��
�k{�]�k�񼲾��	�4'�"~�9g_�;�1iZ$6V2�@(��}dr�4��U����ݡW�29]#>8��%3S��GCݕ`��%�n�Gl��\�e^��|����}� H������Yj&ը��*z�N�;��C 8а3�����M[��C���Yn=�4fy��=y�������ѣGYb��>�APL�=}�L௼���o���,Փ�L�e�ԗ�XN;�¿�t��1��}���l#�**��S8�6ڤ NN�zT�"r��6	TX�J�BA���ˆ��VŴ^��ϙ1�7�LL&�pP��Az�\�D� 	�x������u:mi��@��gP���Zi�5�}��Aj6�Q�*Iwy��|��ד^xaTߊ.]�P����jY\݂y�v6S[����y�}��~x,Ҁ���/�����y�?�|F�bG��q�ؗ�� s����Xz�l��� @���n�$�5�$(�;ĕ��݉>:_=� ���e�m��!W#w��;���,��h0�<�5��FE1䌥�#@?}�:�ó�ꠏ�I����b��TM�̆:{(-�E]#�M:�1E�@N9$��կ��ꟳ��[�!'��5���{�áFt�&�@(F�u����}@��A��,�F}J3?�{��aIԠ]�����|x�={�����G�#�?�= ��~F��!+9�,Y�F<'�l�y��\s\��kK���C�@��9_�k�n�>?;#�3-c��D�����ҳ б���@#v%��� -�, �v>"�bȁ�"����I��s�HcA&��r5���%*]X��hP�*Mд��^��GƦWM*4dWKӲg��d�0�4�U��G����I�"��X�@���P�@�����{ڞ"V�����G��.�$���~�F��������a,q��0�U�'���@d�:�$"2v,ņ��
����15 �V�}���$.��J���1���:%�`��� ˮ~���Wt���֞P��k���3�N��d�3�4-�z��E� ��|E�H�&P�6.+�a�
��ԋ�q�����~�J�z��_�;w��\�O�E8��**��y�sY[[g���W�"+KK���7	t�ڛ���_����L\��?8L��i�Ԕ�F�q�G��~655�@bI?�Wv���/ȗ��e9~��ͽ��!������v������akF2��s:!T��U�*y��B��v:�������?��	d�sz/�t���m]�y��AR�v��n����[iV��Zk�x�0��/0��k#�j*��7~�~筋��F����)��4����� I��0��b��,�I��� Mb`��2���kz��0,��5��84��gX�����P��V�s�FC�V�Q"X�?�\��@��;vG�x<%�Bc��C�3�0@2�S�v9Tj�MG[i/)\?�p#�	�(P	^�s� 
	����b���r��<��4��q�H]7Ld� S��&�ĪR�eՃN�@�d/����74b�ʔ��b�|W�t�r�(��/<!G����M�٣��(�cµW�R'���#g�9������1��MU�.�2��l��Fb��1l�GV�ȡEy��~����Ј/�N�Ow6]/�ƞ1ʅ�p��A:d�	#���(���9{��`tEH��nw$GϜ��5�����'�6v��\U��}V/',#�\�O�|d�8�y�����Sհ�Rh�K�\�3飯|E��4^m�5�e*�r�s��Rf�Qf :w�y@���IN9ϔ\�_�������|�5����1Tpp�(a?�Ҫ�c�~���3��/{�$�y]	���gV�������H�~HQ#����b4����bccgB��s#vcccc���*4C�4%2$͐�HI $H86L[ �}y�>������nr6(�1��bwWee>�}מ{�q��(�C~l1�TTK���0���d���c��! 㬳	|$������Xy����:���{e|b����T�8g c��uX4�hY[���A`�JI'	�V�� **�ʐ�4�E/��������YuB;�d�3�DB���q6੡~���k���<�
ٽk�\�r�t�AT˲��@��apט�;�X�V�
�����f����\#_ ������w���R]����YX�Q!i��3��i&[�`I�%������/���ڃI����!�B��}������������g�}~�/��J;�O��@U����i��фR��k�����;w�����ѣ��=�����6O�ͼ �'ח�&75 Gk��1�-�1�	W�'=u��iл'׍�e�ӞW��[?r��|L�'w��߷LN�\�N4�D�3���|���X׏��=����NC�N���Xb��M%Zp�D�\LW2 G�؄2Hݴ� Tr�bf1�o� Ih�ֳ�!T��Q8�����l�l��(�T��_�x���9r������Jz٦���:�\c'U��E�3ow"�ݰr#��	�V@�vZ]�����;���l����ߍ��V�����])��U�!Ի4;��P~�K�@l(����y�a�t�dѓ�憪X6O@K���n�Ary�B�� �s�r��U p0;5��v7���ںޏ��s���9�u�Z'�c�`�cZy�J$�:�����J�@8FǕJ��gT� G\?#A��i6><6�^7���\<n�C���e��x���jeXv��-K+�tVCCy����<��:����wG�wޑ��Y-n �e�� ����1ٵmB�|Uf����tm��KR� {�ɕ%T��ur��{�(�H�2���- -�Xٚ�+j��YXG�I _�e�'���j�:�n��7F=�Xk��ȁCT8Z���U����MHsU��� ��=��H�Ǎ�ƈ� �����}�6�{>r3�8b���K�>kZ\\��:s|���&�Yf��!�ѣ/�<4� ��*��	`@R�0��:VL���r1(J��f���]����F~`�j��0�Yp�L��"P�[w�Y0�\�y���)���^�KV���hG�C��nM����n��Ҋ��=������,��(V`8� ��gdǧ>"�֚l۾Kz�}��s���1Sl¡��GK�#\��S<�r�M��>�-���&��G۬�w7@�ZMuҸo�?��۴s�<������g��g�������.�,���c6�e D�b=�����/��W����Hע!�Q���~�wd��&1p-}ny�)��^�d#G@�͠gdh��`v���@6�/:ҜȴX�1Nz��0� (����+~�'&L2%N�2T)ʪ���~^��$��-��kPo����=�z�f��XY�ک+3��t��o�Y������ȉ#�IL�az=��H�[�8P��K, h�"�\d�pǔ ������2�B��[���%��[HXg���@�Q�eM��X��m}�?0��붺���Y(��A��) �p����J�Y-��]�^A)���s�|�/�"�~��Ԭz�:N��bGe�rO��`�h@�~?��q<�7��7������7o�O]��95�4�V�	��ؽGq���]����j�#��Al�^bF7���\9wNfnܔ��O��G���zG�'�c��F���bl���E�m�����EbT��?2��'-"w'�����%4��e\����Q���r\,��,~=����׿�y��ɑ����{�9v���=�?�����"��q���U�.��Y����xVJcS̆c�"��Z���$Ь-���"�����FJ�R�����[��E<�{<T� N��b�Ԁ��y [����Y�}��N�U��N���Z �ѻ�{����36;l��F*eV:�پ��$�^��DOʢk�*B�%��џ�q |!�DR�~��G	%���0-�߱��&P1�ݽA�ďj5���8�� �Y D�պ�v���1<�%k��崮�j�����l�2=r}.�|2�u�����8k�!�*��3|�h?� '�,�2�iֿy�㲲ִ��t2���b��������ԑ]�1+��~[��\�74��&������٭����f��������!�ؘ���}#�JZ�`2"ͶM=����qB��	��z��2��>�)�ڴ�S����'Ns���C���ĄbStX����ͳz�wmmM�c�<o �Gt������ATA�`$g�\�\��|u�c��,�C`��efc�ւK��ӹ��;4������{趎yX		�Q�!�W
n��a�`�;���XI��Ja1�W�a�ټ����v��p��%$p:t��ɨ�>�{q㊦8��lhU� �Q��U�I�+A_A0t��SF�%^r6�P&�� ~:�Dw��N��!l3逑�e�BW�����z�So�N vd��9��c2��F��ac�v06��TэRA5}�.��B�� ��T��3+W��bT��i�Ѳ,5��I��n�j��|�����p��6Vu��r�^����*&i���QL��R�]�疗�������nJ�lvlrZ6o�~�'�|��/�12�]�-w�37dyI��v@ _�Z��HE�ܼ*��r����`M4�oF!K�KkKjG��y�R!)Fݗ����\0 ���*�@5�g�òda��Z\	�2jǶ��-d��	�9��Ԧ	f�wi�q��	:�_�ܯ�G����+y��{e���j�rE�4 ��I�R�@L�%��YA�u|x���8jɸ��r�>L{Ҩ�i�s�ED��VZ�|
L�Y,6��G �*$�Gg�ڂ����j�(����z��+�������j,��P1��ĳD ��R��gD��K����_��,΃RwŰ�o��NC\4��2Z����O��u�މ��`�N�r���W��(�>%g`�HW&!z�9�t�t���^-j�q%T�K)I��{ƀlX?9��� d7XC����m�k��2s�::����<�_*#��3��}zG���Gd�����X{xhG����]��U��\�C�:a�:�)�m&��h�m�]\������hUvn݂;������`A�r�������ē̹r*�Y��U"��Q� Ϡ�g�+u]߫˫�����V��<���OL��Q�ʱ'�5H���hs��]�Q8�p`0��:j�7M��}����|F��m�p�jW�jC�/*S����u�z}��Ò_[7OK{}��F�,yL����x��M�}B��{簵��7$9�4��$!i��JMAK���ٵ�	P�V�`�"'݋%��g����MD����wA��g�~�����V�eJӦr���K�:<���+C9?Z�8�(���R��6�2��Ž�?/� K���W��Y}��
�� s�f��Lx%����8��Eq��\�w�Q'�e��.�0��9%��*[�7��3�lA"`|z�D���R��4$0��g�`���p��Whr^6G$p����Z��k_��8��~H}���&���4��"FmZm#rz��$�|.w�����������@����R��DZKݰ��>x����ڠ�l}aN��62�Y=��:�:C+5��X�ʅ&��y���5D�)��p���Q1g>��g�F��l`�u���-��Cv1��Dv	��}��[�Ť �X�P��
Y��4������m����zX._����R��N�I��&%}^�E5�j�+CѬ-[V���}��rD���g
򙱩Ii@�hr��A]�S#�Hl5'
#E�b��?V.�g�Bd�
�n�v�������h!�����.�y�-.̫ᮋ�%������7X��麒���� #/_��<��J��jWVVn1P|���#����gE�J_��M��,ʖ�(M����8�@v�	S>�&�Bף���z]e5�C\�	i�l:�9�X�^�$�����Q��cA�R�5��Ł%�Nu��!�pQߧ��J�(���u���ٹ{8ʹX73��ʺ���Y�$,�C��^���yy��I�����ő#w;A�@t��7���σ�b�W`������@�a�TV�W4�Ѡ�[Kl��!sGkB�t�<VkB�.����W��_���P9#Fr�ð_�LS�cL�(����}�˿�y�|�����ȼ�M�%��������=��\�[��ٯ��!ړ�����
H��^�������o#������=�I�y�nU�&R��X���l�P<�o Aj�I������h-\,�
W��������Bʏ oC��؀�A&59+���1aB]'��'���᎞{�I���8M|Ui�f�dOܖ�-]l�-���l}3�
@��ҎU�5�C/��\$xO�![���x���= ^�Dx��W�vzIG?�Zį�z��O�z��>Y�5������^^zu�"�A��pFn�V��¸�#�*X��E�rD�Xf_�=��͘'D�F�>�j���,ʂ#G9��P�X��|fJo�d�]ӻf�y'�YC�d
Q�.�x#�1Ƙ�:�{���D�f��[��եR�mG�q�3�pM�?���ՠ�j���52��eR���V�	�Q��}uR�tHGZ��z��#J�~�'�D(������q̌�d),�֕���#s����jܑ��A�
��f�*@A	�Rk�����gRIG)�6lxR�ݛ/081�L���p�qH�)y��6U4�)b� $DQ����g������w�H�@q��`��-"�A�z����l:�jп��S
*�m��tS�鄳@/<��.���wW��h�B�J�5]S�T����n��\ �GE�ݨ�:��m��=*{�H�t�>
�S3��u���>�O���a>(q����b��p��87�#��>Q�>>:N��><:"���0
����=<R���Ͼ�*�f����n�Y?*6�^45C<w��k"|��0ܦY/Ʊ�'�F�ILVա�:D��gLMofyn}n�\�F܂ʁ�b�=(�u8�2�[�@���k���Srϑ��/1>|��T�ZϞ;���Р,u6����  ?�7P��c�
d���`o�i��G�	��س�<���2�y3'!FJU�t�|��dfq��+���7��ِn��Z`r���ݎU�����"���(�?�<�W=CE�셋���!b[<�kl�$��X�0?�7&��~F9� �15t�Al��_$ ��h+����fKn^�$�:8���@%�d:������0�w���tvr|�?m-��Z�vC��	�����l���R����(a�Yp�p�Y;q��2�Ͳ��4,q��z�mu�-u�L���`A��G�l�f�8T�	�I�*g����@��I�ӽ�W�S*�"Ki�p#H�)��3����+ �h�5z�=��݉d��\V?$�8;��+�f.[xshb����^�i\�{�Ѓ`O��_}i����k[������F���'��0��q�.�ڶY ����P�]�A9ZtZ�I���}0d� x��+�|8y�Sc�BD���)[Y`���$'�d�ےU}�ȌكuJ7O���; QE��Ճ�#�;1�
�O&��ɚn ���C�/�yE�u��4�w��# ���LAN��6��!�2��NAf N��#c.+g�*k $��{F���Cb���L��q��
�*7{�޲ bx�(�z�E:�
�KG4{s�3��b[ ��co�!��'���0X�l�{�DP�*g��(tR����2s٢T��s����
�WKT�m��ʪ�]SbWx��Sc�rϓ�ɓ�?*{wn�3�~�����kD��g $��� ����P���C��\��K/q%z���씫��h��bc�Rǃ��,vfC	͗���~����82�,:8�y{�1˞�2KL�%<��"~�k��Y5	bӀ��9==){vo7�8u�#z�������:��~���
��vc�N�F�`��r��  0_�;ΥCf�U���`v;��B��cG�!�7:�P=
�����d��+��~��}Cѓ����~�A~��a�1�k@1\ˍ��U���!��

�>�@����郶�2S7�����c�6���s�ݜ^A�����$$�c\���c�f�ʑ���B`��:�"��
������ �oM����M7D�| � ����6�&�L�A'�;��ĕ�7���t��ڲ����sx����ɓ\B����ݩ9�Zc`$N�UG�Ϭ�@�gs%�}�Nd��B����>pt��wMn?9;;�����68���箁N��'P۔.-,�����|���ϟ�&�n���_���
p.���7�ާ�߳ׯY��r��
���WW�z�?���kl׏;�3��P'.Dќ�B���nԌFoЩn���3Dméیm�V\�^Ǥ/յ0!xa(,r�JY�%+K�,�&x�����(��F��]	����.��H%�T�j���~�Ȫ��A�:�P3�+TV�*ަ�z�eu~7�j��X!��.Vh\�4�ZWA?YSU
͚��R*QjX7��͞�,-�鳗�Q奡YGi�j�Y��j��&���
���B�5�e���$%��pyĺ8�/Y��?�p�?��l��7<6l�W5Cyf���%��f;�.]���}@�:x��?�`���4��{催jF���0Hn hVج�Q�J)��#��Č��@0S�v{���=mk�C��N�^�̢G�/K�F������>);�LQY��F�ѻ�˓�'���K���7fg�¥�jP��ȡòk�vW�<==Mc��/�;:v=���Y�s�X�^G΢y�+�Y��j��M�>���{���+�Ȑ���%�:đ�{=��^���POt�gI���$�[�[����z�D,�����7��=:���K_�VqZ�����Q�� K�g��J\���gr���d�����k����ޜ����8�Rh�sp�tC��a�S�D��h����wVNG%���u{��������7NH�Փ#�2�,�����2�Y%��n^�*���1޶��B� ���"�'����՜��i�4�߻O�w�,X ��q��|U������˯J���=d�	�!Y �
a���<�,���t� ��-h�S��ܷ{��o�ݜ�*����`��\(J[�,���Y�Ե9���2�Z��9�M񙺓G7�S7F֌B��O�vv��X�s�ޯK�zô& }�FT0�`|�{�2!N\,2Y�{"0٪�H����O.���oq8��3#�	naE��s�g��u�Jut�D��<��B�eY��8o{6�`S���!�{bF3��]��<�y\ȓ�� q,y����lR��i�^4��i=_�uBu�QO]Y
5�\�P�/K�z�T�
�BC�:V{�X\.��Ns���ϯ�<|���O֛�	l�Qu�C9~�M��)��TKe���R��͸g�6i�.q�d�Zb�;�%>55��IY��V��~�{/I���"��}èY�(CY�e�ӓ(H8��1�G����(WF4���1E�C�Q}�!�jhv~��;�O�����:8 �Nbd���NA���Ǐ�f�X�����ʒ~����x�u��0�tcn�����e��1�jp3���G�����'�଴��M&�#���Hq����o� �uU��~����Sy�ߓɑ����*��}��oݾ�����%��_����NM��}�)���?��_S�F����2��օa7 ��=D[���|���Y�q�ߪ�;XZ��˨8|�}x䝻�i���ߛ�4!O<��%ͬ� �B%�\�ӡW5���큮�,]?��U���F��Cx�{�e�vcF�zo��b���Bdzb�������+����^9�U�����7g��k���{
Q��ڼ?&V���*4���Pq�B/9_���?�I�Ϗ9@-
Q��R[J���E]'�9t���Oex\������qyI����Ѷ!��e�i25^|���y����{�%gTp�@��颼|��yy�����oJO�kp��`L����NM�%�D�@�R�%2s�,T5�$�&5�<�=|��]�?dUq۶���c���GǊ�F��C>84@[ ���`��� s���qC~��u�u� �a�d�u�/^��9A�T(I��+g��I�}��������.����_>�3�>|�ѥ��'�q���tڽ=�hUF�<�����g#s�&�rJX0��El��n�<�ƚ.�2	d�_�&�7���i:;D��c̨`YH!�a_N��y�|���g_��r�
A���@#����5h�
Ia���E��FE[�ݗ/G����Ʊz��ͩ��s�o_�y����2�����
PU�Ѹ�k����H����Nk��+V���)e�H�~W+,WG���N�F����w��;���Yi��P�:1��h��Ů�30��O�sܼ�p��pd�r�W�!!�Y�{����܂�޼)W�_d&D�}�yu���J�q����h�ڙS�����^F�0Wy�ԩ>(����e��U��j ��~�Ta	��Y5�h�#SFI��N�:��Ϟ���J�~�ƮOL�����2�ڹs�,޼J��RN�U��5�z�dێ�쭧�/�?�ň�a�tPnͰ��G0�kgsω)���fhD���r��a��t��{��͒eN��f����1���@�z��Z��L��1�=o�}5�gT�z����5 $D�F���g�%��&Q�֭�Y�]_�g�CU� �߻`-��4pC  �J�V ��������*z�~鳟g�<�5��n��:���fϺO�ڷ� 8ɿ���%�՚����,�#�F�U]o)�qϔ�29����^~��  >	��PBG`��m����,.-�u�h�D����l٪AC�"{v�auS
~����&�Bl�`H������v��G�^�3@�ib\�ٚ�z�<��eI�w;	����GL5���o�q[��7y�������}� ���2�	�3�+�UӋ��pO��9��4x�X�ޯ�>��gD?~T���e~g|��c ��}��c0 �>>�%(���{aH�h'�4?�=*����
ۙ�P&�͝�]=�Sr�m�w��t��K��u)�����Pn.�f��S(TL�8ut���E��K)AH�Q�H~e�6G�v��q��#�	؈:J.�����OL�O���x�����ſmo�E�뺐ko��4���ɚdb�\�m�|`�`@����r��=4kh�$�}�Z���"(�q��¹����Ͽ"Wf���Bƴ�� �������1'k�S�U9���Y���ҿcy�="i�DQDg_Z�������5u����<g�evnNN�<��G�%u�I��7��`��&]f�^rR�#�k�{d�7o�\��^�˗����~D9@�ȴf���a+���vD�"ќX �T�hl{(k@7^-��ðep��!��$���� $Fguy�ƭB���	��Ƽ�Lƍ�1�enU�`��2�'��D���`7�3��D�L~���HѠ�I��5��e�Y#�k�@G ri6�Y[�����n ��w�  �Rn�kv7,�ϝ�u���Vz�'��jAl��ݷw�l�ޢ���)�!�[�
�43.�I�E���1
��zbţH�e�F\���/�r�o�����[D0!G��i�k�i ���\[g/]W��A�]r`�nNA�87�%z>Ș�቉I��3�ն��5m�3�,Z��~I��^��Io������)9~�-�ݘ��!J�-��.��������
hw�ځ!b�j#Q$z�kZ���׏������F����:��>�����F&�A�����
�Q�3_5����B��A����'HIM!��'�A�Fbp��J$�!Ԍ@VG�+�S
��9���=u蕇�����/���+�כ���^�)f��٬��n<ƀX��2�zc���F	�X$�6^�԰Q, $d��͹i�t%��|��lid��������c����׽F݌��n�B����0��7Kq��꘷֠�} �fհ,�������C�����r��U�]�0��.k�95d�f���L����m���(���Z+P��+��Q61��w��.����U��q�ojF~��uVM������\RC���P� �,3Ք8� �yKB�oanQ^�l	��Q'�iv����6���ϨTJ��a@6�vs���Ŭ1��������3 ef���uB�{�9ٽuRvo���:7��"u���^�:#��}ZV̒��V�ߜ�#w�� ���r���>�yƕ,ayX�菠e�}D�OO��0Z�k�`��A�~MeY=v�A�'��~�A�w�8��^{�u�K�~��s���A�.�^��1C#�7��=@	������~ܠa���,^�K����p�n�o~n�Ncxt��m[Չ�Hmm�Y=��5k���p�)NW2��-55E��zO��d��[f�"E �8F�0� )@ֿ���0�@�1vњ��y��@�����C��[6k�Q�Gc#|˺N.҃����t,x�;(����SGϞ�b��@e����;�Tpۀ� E�;U�3�T9v�v8it�y��Y�û$6.�)�]T?����r�*m����I!	�c���q	`䡄�F����C�l�U�:���g@9��Vtt���v���H�2��,��d!�޹Qeh�Ʀ������;��w�x���v�9�R������ߍ��(��s����&� �L��3�,Ǚ"��CgH1��u�)cL&O`Z�9/��hC�Ε\6���P�k���]}7��s�`�@ ��K7~�����t@]�$�1>`dk��O����<�R��E�Hu�mu�m��t3D뢽 ے�42"��f�=J�N�=�q��%n\���=`/@�N%B8�K�����������������[2�9r�>a�V�٣G:��FX���9��|�:���A���zya���M�����zny5� &2��y���2�ҥf<�t�A��1�0O�� �n��e�����<sZ��]��L�V�clp��F��B���#w逳�����sT���+5�]�yϝ}��� ���F�=p~4�ޡ���-b�/����#]��	�H�2g|��1nd��o2���;@R,�n�� ��gc�ע:�y�X��������[�N:�W۵|6�K��ߨ��|�-���g�c&ȭ3�aPZ�{��\T�@|��kA�ڂ|&�f�s,���G�C'�N��}�:X0��9i4{�B_�.��aj&� ���ֹ�r��u�]���ֵ;���('$b��Jz���J]�t	m�UK�nO�=Oє+׮���
[�1����C���րEa�
����"�q�&H��"v�%n*njd�����6�`> ��S�f��k�C&7Q��5��a�vy�gb)�0��en	gx6n�V�1"������tmU�0��&�S�[��n�(����C���ܡ?�L�����
��͛�}'���{�3����=A4�,�J����8ǒv̞�v�z�=e��8g���,���k�P.����Y�ζ}G�g��(��詳��Zo��'F�
�.('��i�%H���߃66���742��S�B3�h{�)��XD���:�u�zY��N";�L`�'ވ{�
�s��]T�	@%p����tJ�lx|R�',�20Ʒ0�#V�hӥe5����	ئ�Z�����5�L�J�S�J4��xf,���9�J�(t0�ݓ/��X���ڽ[�t]����u�b5�N�z�ҳ���f4C�Fk���={�oQ*F� 2�s�E�w{��4�C��V/��F&y���ߝ�� �� ˛�!�٥G��L�#�}	�n�Ko0��7��!�i�yF��`w�{��|���L6
zcn����>mAy"f�Md�0�Ⱥ���Q���d
��w�u�\��� �,���tb��e��&�:�y��j���F�7[b\ ���B����l�C�y��)�r�����~��t��8����$&.���.������/��R�>�Lq�����p�K+�M�J���,��������B/"N3R� uyy�{cd�̪�{U�l�T{�+N��4sTI�����@Ϛ�\���}��L�qPb�>@,?���q��A�eemE�&F���曼%�V�?V�둬g���A��ۃH�~�F]��1�C��gW,x��b�F[qѡ+�#80Z�;%�w��{�W��������f�s��o���#�o��sA��aJM5{�~Qa�1�����0�+d-�v��_�d�K���8���o��Ol�w��n^�D��̄A��)�}��o����@���-��}�����!(�����jT��s�f]�6"jl88�MSjlF�IWj������yne��D"1ptpxW�
����'>!�G�~�oԞ#Ձ�s[Ď1�5��i����=r��E9q�����cg ĩ��عC>��ԈOW��e@R� �u�T�i��UPb����D608[�78n��$4� fM�W$�D�����-���tF��T�Fnue���Y����s�I�TK'� ��C��U��^k<�4�	��eh���p�a��d�d��,�(�:`��p��A68o0=���A���O�s҉s�D�9&aV��g�'΁����6���I��&�o�������=�+n��כ�Z�{�Y���o
 7������9���{�ʊf��_S֡���^��jI��18k�~�������bo���G'���Lph�Zu�!{�墁�8Ӯ���CK`�%8q�u8i0���u�]���k]WhW�� 9V��C���*��rP��=)����lf��}���� `j18��LB:M@(1�)o���9;7����X
�z �a�C���2�9C�c�όt7�P��DRI:@'-}�b��Z�=#<��4j��z�Q�?���\�x�/K��V����^��Dc��O����^��e���=}����o:���vwe���Z���|�H'�!�m$�Yc�"��z�a�����=��D�\�lo53s��^���b>W8W�K<��^�>�놺�@Z�~D#|5T����m���3`$��-�2�f5ȨF	��Ҧ&W.R��"��O�@���7ݠl�����dV�Ҟ#h :i�"M5���iO�n��۞ 2�h�V.�4r�JH��3��(S��u:r�o�����+?<&75Ӂ|#�	�K���,+[�얧���eL�5\hKI�h��^Y3%:����P�,����1�L�j\���'�$#Y��m%Z��D�< T;`@T)rD���Q8�L��zju���2`�]������)���u������'�tl�,��qx&4D����E� ��L<���Y�`s�d}��G�GLJV�ښ�~
��z�aV�����J�sh��կHd��>@��<�gԙ������rUj���7N�$�{��M����-�ᡢ��sϜ;'ud��\� �XG0���hC9	�`Ȧ����6��|��&~baa��javN^y�e��{�aٶe;Dd�p��Jx����?xA>��ϒ��l�i 3:6L�?��/[�/�����G7Q���m�w�3�ee�g�~�����}�㟸O��w�<��G�����{���2⌷�)�C����#�I��R�Fȃ�F{3���B������5F�����4��^�MV%^!o�A�A�?NZ����Z�_V���>ٳo�\���ՅEVOP�A`�	�W@�~a��.�"�s����k��P���s箵�����kwwZ���ApwE�4h��b�X�Ȫ��Aƴ���[������ޙ\)wLM��lv�f�X\�{�h��<�\E]3f��I'��:1c?ju��!�DI1'�����g&Cj� ��jf2T2҇����,n�iQk�#.���#��4"i�SUc��Yy�it��5a9V�d�^�nA�͕yW�;�=�~9�`�M;��ω�<F���lbF\�J���QU�
Y�lgU�{�W�����W�=�L.eߏB2���8`
�S(�}*��35=��]ZU�>��L:��t�= >���0p�!�IȟM�� K��G���\PC
����s���%#s�����3�WMC�ה��r�7Ͻ�q��A��o�ӣ�}6�ǌ�ԟD���{ �'�&��mC�)��C��X��h%q�կ^*��a���CƖ�6�r�%:'T2��Q����瞓��\�x>plk�:ecyh�@Oh��]T�戚X6���J(
�gp}�z�J��,+E���?"����D��F�^�d߮�6���cyaV��{����2i\C�Z�����xC����/�����?|T~��klp�"_��y�=t�fUG��{�	����� Z��9z�T4����2���ΐ�{�h�0π��������Ι�dyi���VT�̡�Pl�,�ہ�2`�d���-s�eM�2�1+MX������)���_s�_S �zѕ�|�� �w⃳�}x��c�������c���(f2���`�	��mR�̗�顿��Ϥ�8 ��K�Z;u��\&���ݜc�^4�M�_�2P/q]D���,�EY*$�����_�����G���rp�l�g_;!'�zKr��.��t�I`2o�c|
Yz^��֩i��C���S�Pzj(Q�Ix&�nuU��5#��F���Y%AcT��б�����8����Ͽ�����6���i��,?ic9�7�lb�2ipA��*G5�(s�䪻unyM�x무�!D�q��c�C��J�uuiM~�_����#c2�����~� ��\��^�# SpD6�]�נ-g����$����A�d>K���4Ç�K���e��+5B
l���ɱ	Y[���ù��5^��WN(�jU�h�	AyP�yy��r&�+���{�Q�����Uڠ��`�dn���6xp`poY w�3�P������a��H�<���C$9���:
��Y����%P�&Pl��&M5�� n~iY2劌n�"�~���$��񱒒ϑU�o��R��<�>��Bi�س�m��}+����ϓ������ګ�p4�c��l޺I��e��7�"o�;��AF�{�e�V��G>&Ց!�������޵�A,�'�9�����'� ��x���pߠY:��jk+,-��?��2\�˿�7_���Y"����*y�)�t����˽���ٳ��O��g����r�����o���IΖ_�r��� k|���<ih#f����Q�s\׀�pʤ������F�躂m(dK{k�B[�(b���r͠�R|^�@�5���V�j� �� t=���%�=�F��|��` UKhd�j�1z��I�R�1D ^������g��9ztY�X��N��rz
�+���I<�3���ind<�t�������K���H^3��I���&��F�mS|C	���{���(}ayYN�?'�φ�v4I���SB")4bh���B~��ʺ67=4Ta�P������u5C��l�����,^��Q1��46���!1�jӃ�B_�Uc7tt���4��Ll�]6�CA�:59%���rsNFA���'=N�q���g�e��u�-���EY���~[��j�Fo`���q���҉���b3ڕ�0��g���`b|�z^�,�)�cZ]n�X
��)A:Ru�� `-�$�VJ���僙�G�))x�^�˟�e�A���*u #�p�� �2��h�}��1= �����I�tc���!��nA�euFH�2Ku1���]�%(��}T��9R\G3h8�}AV��3:PT�v���^5�ѱ.R��sI+zm��y���"��.�v��߸q]~��O�^���̑�e��M,+�9s�#� HBMn��W��ӟ��P�ݑy8�_�����=<<��9����E���C����� o�e��׳}��ܸ�(?������2�ܷk����C��y��5f�����o}�k$�0~�~�J�]�������Uq����$���[�&�҈�w��H�m�:�z�p�3�]����y��~Bn޸F�"�OP;�� �_t+�s7���/�E0*�V�L���Y�Z��	��5>������u��Q� �=8~����g��KGS3�z��6F���ݮ�iK7gB���I��Ш�@�A���{�T6�}��4��9]䔎,�&4� ��6����_˱�	����PH�"F����V����f	����0�@��A�9��#JY���H!ň�1zv��@�kf��F��좼z�{���73��F�����cz��H�udt.����ܪ��`w$N|g���H���o�/�"�k�ZpT@�<��^kQӛ�;�0�}��;r����ܹ��i|l�4�˩��AB��H8M �80�M����^�G�&�DN����m���#�h���6؋�ڏ���r���0�M�"a��kF7�[@k���&@��:N�"A+�怅ӛ�Rh&�?_[]��,�_�w��6�?ձ���&��|�26�U��� � �WãU�'b�I�ʐ,.��Y�.��~Mf�_�@huVT���@��A�!����;�_����"I!]�7@�����3-Sɇ���|��!�������,��Ȥ�߮���H��V��	�9�i��y��Y��`@����Qi �.`���B������m�S�I��C'Lȩ)d���f���3��4�5�w0�Y@e@ZdӰ��R���wȪ���I��9&DPA�9� �>��n;��7X�P�Z`^V.��`���;�����\i��Uo�8��2AѬ�na~�z���'Ū�E�u�V�������a�������ߏ;7�'<��0 N��љ�qZǁCS(E����A���QC��Gf���`��<М������gx@�����9s��ٵ�1����4�a$&����=,x�y��{�5c���Q%S=���TϊY��,�!�Q���h�yt'F�Ԉ���I�83//�2�9������_�'�&Y���$ /�1��3��Z5N|G��r��L��s�v8�s����i�DӘѠ����5s< ��?������������}��׮��)�����A�P����j��|��Jd��wԃ�G���w���`	���9w_�'�v�����a�=3'�G>��B�7T:F���V�*=[�'�����;婧��d��ڪ,j���g�#��r�*z^ם�2i�Ȅ�''�����ݹc��7zr��)�?�C�WXQAK�֨�i!Csߎ�i�:9)��$��\-x�@���dA���R��-�"ǖd ��0���3�kE1�j�I�|��=��G�c}��a���L�!�5p��D��u��k�{߃�/��gm=�y�����(gN��z��F4軦�	�����u�u�=k�8��!+y��c�����B�1����_������1��s���z��x�P�k"((�7��m�ֳߕ�37�N���S}r����p��>F}��I>˷�|y�sNe�������ܬ4ke����@��˗� }2��2��!��	S{X�;ǻz�q�?��@_���؜hd�B�dy�$P+���)�(SS��03�ߥ����xK�m������%tD��*�O����4S8�f�5%9r�.��_�y٥�or��YK��lX@Ve�[�#�cQ>�pŘ4���͗���qn��hs��9�L,+�U�J�N8�'^d&�ר�R��*��	2��`R���8��!��*��@��3h�N��0��lrF��ﶚR���Y(���^�u4(��n�CG��c���1ҹs猻@�� '&i��O��سW��efn�._��|�;6h�_~$C�1H��/O:���� �9���Y��ٹn|@161*G��)����@��@iU�D�,n޺U��U�� 8�����\'X e2�;��0���5N0  @���#��'z��N����
�aj���8��
��$��0 �EF\�	�`�@8�s��q��y2�%�-*�(���g�;7���繴&����+#�¼��qA�>95%; �+�����ΫE#/^CO���"�	k��\�|V��� {A�/(�7����;2�0/+�`~(�KW.�}z��/.[{	�&�,�"�{̍��3YQ��X��Y�-�jK©%�s���C�����[����@	{
�����|�S�b������j����E�]��0彀��V�d��V�G ��8�y�������&�f\9lu�J�'�zD�uu��ۜ։9�L�k����N��n��?��q��-�5�#B��.r΂� Ҡd�*X�����Jք\f$�X�LJ]:1�v���~�t�s��&���"nx�j��I5C�)P�+��ۧN����Q�����,�,��vȗ�v��1yJ���^�8�>'����⢼r�5��A�
��D��1�2N�8-_�����1�A�Y�8^��mw:�@Y��5�j�m��:��yzJ����Y���ߡ����P�5F��=�V���#�{����$���䑇�j�~̎�S4z@�nҌ��_�:9s�O?�Af��r���[��,ö2��17���}�����,���Y�����cj��~�<;���>&G����+W9�g�ʐ����۳���׮]c�NY4�Sc�t�����{x�`/��!i�><s�'2�N�+�(_|��lQ`� ���i�Y�b�Dz:��PG�Rw��R�k8�EY'���wŪq4��N/�����o\9�`j�u����5S�ӿ�ŗ��_%�������V'�A��9mW1�H��CD��1�O�Ξ���/	x����e,�*m��4;�- �������u��|�Hw\*Hj�ZbP��k ��� �D����;%^{�\����7��k�˿�Y��Q�ܔ��n]���#o������r�����2�ǔC��An>��'�)��=�dm���3p_1�}���`�hp��u��IB٨!��i�%���;��$�juJr�xW�;�'<J���22�+m�A���l#J/�\�c�k�9e:�˯:C_j"�%k}dO��L��*�9�`�I�����L`$2t݈>���g	�Tq�,�9.G|�կ~Ք�rF�Yk�C�|���������P�#��@G�{vq�8�Ӯ�j�
jku"g�*ef2���@�l��5!jA��4��	���;x���&,	�Ǆ�DD@�	��zHFG�\}�q���l�
��v���k�q���ٌ:k5�7�\�#����߼��ڕ�e�D�s�=�q�M�D�"�x�}���n�;C��Fi��}�h8i`�{:t��{ָ�``p����s���&�dj��:`�mS˞������,Q��y�����Q�������lX�Y1���zK�����-�Kn������vA�k k�@?`74�o��E���l޾����W.^"���9w�#o�.1��ۃ��٘aЃ>(��������g�^�2i4q��#r��!���"��������*g������4���J��N�;p�Q��4��꒾�E*YaЎ9��w����/ʙS�eX������,����%޻�z,�~�C��#"����I�{Y��H�U+
���M�f<� C!�W�\��-`�� 4$�{���%nSRt̃I���q_��PY�s�f��9u��~��v�WOK�+Kޙ�Y/�k���ϟ�(�4�3C�*��٘g7�Jgr�.w�OxdK�$S(�kS#U��%���Q8uz�����l��&E7�J�e �@�O�gjb��b�ǲ�>#,�dT�#a_,eeV ѫ���������ₜ~�-�g��a�� * g!���jnw����6,�p�$�Q#S��4�	ho1�����h�d5]�W�وJ�y������xht�0!"����M�%u����E�k[�4��D2���*�,#�46(��Ɖ�R_�g/+�>|vUƞ\��⽶��%��}?$�ܐʚɶ�*h��w�f��>{���ݠA������}���~Сߎ.t�fd��Nz~���7ҝr��]19ZD�#��P��`eA{�<��;<2*3�sԺ�\�@�����K��}F�����=��^7�A�� �[A�p�p�4�ff���YL�z��)�s���@v��'�\�UP����'��?<�����������^�u�����6�������?��_'�@W1&���kP����IW2�d��fÉ�C44+ַ��܅�.��T�*	d����/Y~�Y>�ɏ�3��pľ��o���gx����z�|�WŲ�bYr�ܜ�б��*�-p�Bɥ���9�$qІ,{����c�6�y5��:+b�:|�L躽z�&�%�3in#��G���b~�Q�����5J퀁��_���^[��l��o�}b��OqLc���0f��0L-HS���*�� Ӓ;ǻz�q�?����^��5���z��۴�f��Ee:��/q��x=�W��ID�gT��N|?�>�M�HR�Ӯ��gO��o�y��X ���/�8@ ���G�(�M��$ɖKd]�{c�7b�@�]Qӿ�H��c�~��^G�;+�L��u�1߮�]d* �U&&�0l� ��qN#geu� �q֖�gm"�1�D��!}�qA�9ʞ�]P�����^�!�{vn�Y͖�|�S�g70.�0Mw���{�����3�ȑ����>���i����� j��)t�@b�Tv�<&�F��,����N��-��>�2��n���o>C��ߗF�����|E�Oo�׊����!��A�g��s��9+Cx>�~S�����{5�\�o=��,,/�u`�s܉㧤��������9p�X�3����O���������|2�U5��������p�QAB�sߑ+n�>|�F.u�>��ﰕu����T�V��~��5�v��tm]�x�����y_���y�;�bϾ�X�<~�=����_~� �s��<�I�\�?Z5���ޛ�}��R���#�Y(eI���˯����/��\<w���5 .5������EH�<>V"�HJ�<0���z ��^�q�^���U�u{����y��{� ���(��3�Q x^���A�`*�E����>�Ժ��?G��}<�R'���MyVـHU/�A��̪��>��[���e������C�	������R2G��dG�xAl�.��C�D�n��<�|�a���8�,n\�ɹ�nd�1q�}�挱{�8V���=|�@��_βǂ �эƠ"�IR��k|rDZ��V+T[ۿ{3#T0��e�4G@@�k�56:A��Z�A��@�P�ڳg��(�ӡ놾r�AX��E_��5�:�;	L�,:d����z�4\/`p=E �H�ˈf��>� �{�獲.z���L�3 �gp��U�r����55;��WY�?x�`_�j�������Gz����{��c�v{��>��ǭ}t�㞛��� bt���XJ���"���_�����S+k@U�댾�9`E�8<`��l3Ḧ́	��xр��wueMN��ڶu�����|������ҁuW�VA�c@�6U�PeIm0w�I�7�0� ���/}�OeP��iէ~?�Z>�����S2� ��AO����{}`]���8���r�E�'r���ݶE��d��Y�Ԭ�ę�"�D�Q5뢕�'ޔkg�hF�c��P�`~C[leaV����p�{�2���\8T�b`���=�Ԉ24�[Ce��O��O�>��Jڡ�'���+�:Z��}��S�o|���K��#��q21�� �h5�d��7H��뾚�R</�2J�:�������7D�r}ؓĩ�e#�&�:������vg2R�!5#����.wn�Ox�6�)T�����Nj�l,�2JT4.��f��A,ċ����~*J��#���[ѭn�͏qQ�ȕ�B���"�pw��>At0�������a�*V8���IV��`�����?�if� ���7d��ݲ}�N��~��#M����Y���U���C#�j�F���:�	u�Ȑ��$s��eद��{�n��adh�<���~����҆��5u��U�U�w�l�&Kg
���E�Qb�g�Ԭ��
8�c���7ԡg���)�s����,�`����P)
������s�p<v2�m��N�r;˛?n���v"_��}�>�o��J��E`�=q�X0u`�C��Sk�cm�lT��,�QH��R��	�Qk���]+���Ժ��o�;���G)$�
icc������������F|=�l� ��� t���{� f�ggo��W����3�<���#R-��UD�BO��BR ���,����ٲ�?|�u���ߕ���ř+�X���	��T��#������wI���:�/TY"��Z�Fʔ�q���ܑ�5�5p4��ί��3o�w���4۱��*Y��c ��D�QC���ڒ\9�� ���_�b�* fҊ^�9Hb��@���C8���뽟�}6^�*igmtIV�(ṢjB_a������`�$��|d�T���e#�ȁ&�(Hg��8@uI�k릩��/�8��'����9~��C�	����a��}_1a���:t�f��׭^(1�%�bΫ�AN��:��,]O���f�a��l/���|Έ�g��-�ǎb���B5�����> [6Miƕ���ܼ]&�7�Z��{���Y_�'yP����pӮ:E �ӘAH�	I`���fM
�ш쇆ʔ��`��COr#?������R���I9z��|���޻K�m�V��Ȏ�ۙA���PΟ{�}_��#�QB���L�5`�U56Фo���:]D�,B-����@?��엖�4p�3K�6$P�J�z��J�n�����oj���+r�$R��l�?�p�����`p0��� `�s��Z,��W�c�6_(�9�^��Ib<��flݖ�e@d���x����RRַA �De	�s���8!֐fo���|�ߔk�.9�HQ�|�Iy�G��_��x�c�d�K�E�s���\\WGO��t�Q�Y_]d0�B$u@G����_hp:!�r�Ae�����ZHXF���zM�JV�!>E��t��WF䇯S��&W/�����7���u9�g������UO�P�oB8��϶��D���h���_B�O�eD�JC��������r��E2���$y�F�65�����O�_vl�JfC��$?�i3��WN��?�җ�x�.�;�,���xem]���dSw��_[~T�/�oݺU���YM����{H"��{
c��R�5�2���$��	Y�C��k�#�B�l�C�̎驱Ɲ�ڗk��0�s�٠�#�.�QWm�	�\;�8��0�僜�3�ٓL���M�0
�����f3����H�mC�^6��q.ҟҢ�^�t���C�3�&��
H��;�8��iW��2=͙܄a�Cڹ\X1}9�x];�T�L7�F��&5�l6��kTg�lC���P�aiq����J\�C�	��b��r]�	�e���)�8#s�X	ؤ�
��9���:"]<�����a�%rk��:#/�[K���`�����D
t�Y��1q��1=���ݱKFFJ�yrL�6m���M�2�6�����,G�>�ѧl!''߸ WΞ�;h�cc�6q�����U#�]�q��#c�;tP���3��c/�$�c9�i��}˔f\C9�<>�ϯ��O����D���b!�Y�)�Ŭ�!t�3	S�됉�0���uZ�]�|�}\4��r�L=��$�(c�IuJ�3d����ac�0���7|=X6�#@��x��`?��3�ۏ>P)��]�'|���.8�2s�8FF3�X
A���IX��m���jG�������8E���)&�i�ֱ��������% �۶y�ͪ��oA�{@N�} 9�?4��@��P�L/!�1�PN`� Ԧ��ȃ����?��l���۲���:�ߡ��)�D����D����6�*�j"��e�^�B�k0z�PS�^�A�(�q[���o=�:¥�҅*B:|w40�2�JZI����0���ޣ�oR�9{�dS���%J�B�t�@���>��������1��
�h8�@��K3�Ə�`AF7C�\�f�%���������W`���� �+B��������+G�%���X^3==%[6Oʪf�+�Ȭ���-d��`JL��b3�l�T����dr������^BTteUu/b��D�������r�0�6!��E*�4��ǳb�΄ag��S�n7�S�\	�+��A��GL��6�)�?�~f�M��]�ˇ���?�y`f�Sf��XO������Gc	��Y�7[�iL�F�E3�C��_G/��L!���c���=?|A�����A\��a�~�{(;���#"�-[��!��F��(�1ջmY�HpY����:�$��ax��lb�9��ga?�&������%3�C��gܽ*q_�jW')�h(%���H�@9�)�p"f]��}j�N�<:�ѥPm]��UWG�鏮�Dm�l�����a���"�˲}|Dvo�&�Ɛfsv��l2����y�����pEraJ4r}uI
��c�Y���&2Ρ[�������1�}��]��a\3z�ih�$ht#v&PO_�*Cu9d��~i�2hT�]Ӓ&S�V���`�fĩ}m��>X:���>X�����pxP���3���y'�R���g�F�X
d6A���
O��A�����_6�q����Q�hW��P�6���t&���j-f}�4��`׎�S�8���"�O�<���0^�<������?�uC����i�e�U%��t�w�r+3k�%Qh@C	$�4AZe�,d������?�?v8��F��2 ԭ �T)��\YY�Y9o��x&ﵾ��w3�'8ێ�����2o�w�s�����k�	C�|��%��4>x��+��� ���� �K���^���Dl�JBP��j�z-�pZ���{��K�ȵ�����ӫo����v�#g_?+���~_z�A�͙���v��Q���F��A�5Y'G'VB�`5�z]���w�>�ģ��s<��F�ͤ�����i�s��p�RR(|�����)���5�?�<��|����6}K��K�벭�LCw=�I!�%����=S?[]m�)5�F�8ڮT��g�ȝ�`�?�U����/��Y�A �S��p�p(��0�:g�0u�JL�D7�!/]d�y�;���'��E����l�(;�38�mO�U�a|zz��-�Of@'�I&�vu�X���v}�U��N�I~2]�K�>%�S��qS����8x���l�3��O�*�C��&��Ȥ��$���.|Le�5��l���8KRNF=����!�&�2��-�_�2(��JnU<�խ�ac�f��t�ӟs�4����=s�z@�����t�(u���ܑ\F���rC��6	? ơgy}u�Ca>�>��ޔ��ei�!�� ��:�s\��l��>�!�{�0BZV�~C�N\J�XP'��LDŌvp(�\���}r& 2F�	"�2��~.E���꒩Se=D~p��qp��-.P����8����s�CWO��
��y�e�Ծ��xu�'l��F�zޯ�M{�p�!4��>�:^>�j��dJ�E�k���f����)��G[%z�����<x��P�Z9șmԻ1�7���!#X���}�硔�A�"rH��A"w@��9�gN�.k+jg������^���k����h^��%r�demC�ַYχ�QDMÇ�>��c�K�����V����>��<����2�H��L(3��`t�0��=
r�k�t�h�� �p����9
�r��%����C:��LA��b�
ty���p�΁Щ��He�*6�H��_�}�Q�9���8i6}����7Z��tXXX�������G�7���q����~T��o�i=O00i.
�3뽮��TA��kC�X�)�N߽�Hd�Ƶ�%�Uk�2�x߽��^IƎy����	�S��vÎJ��d�t�qi��Y���}�ւ��	+����S6Axk`S�Ic5�2���X������;��U�k�	�@��֭�@)�[��1�n�����`W��k�7q@8q��5�k��6��6܇3��1�H�dMb!j�`����ܥ-j��A����lu��_~�9w�7���KRo�$��Lc��JJ߻	#>��Vb3xr:�oY�=̼puzȤ"�T�-G���:'Ya�D��w �^A!G��C�D`���F*d��|���O��7Μc-��}��iT��z���gK�;my��S�o}�CaVo^�(D�톌4ڞW��'@[�}3�@.�KV��Z4���"ǹ���e7Zap�|�����a�� :0�C��{���g�~��ޓ�"��m�y8C 4@˿�3U�2�u��q�A��&l:�Z�jOVQy�y9�������Ɉz�yU=������J#�Q��羛�w�3�|Z|�4����ͻ6B��|���ӵ�Î~d� ���(T������K��):P��ۿ)���s.횹� �A����#��C��ʲ̶;|��5��SO=%/�����i��F��ޡ��/|��}��|�k_������V�)t(B�/����G��O����/~Q.�}�D��~�{���ID��(%���^(@����3�J�[�֮S��I����Htkk����-�q�v�6���l�Ȧ�V�9 �!E�^�:�GO�/J'�8�����j><4$�ӏ	v����%�k �?�����S��~��N�D�3�a03�lom0#��(�WҒ�x�ǝ��@��"��`W�e�J׽�3Y*����=<����] pt}<�6�+�&FND��.$��%��-�f|�M�I��d�$�rf_/�#":87x�K0�i�GeA�+/�MFe����8ܯ�dC�yy�����3Ap��W�:3��q�rI��.�|I��d��f���o=H7�!v����k`l�A�O77��}��2�&�b#HX�e��ԍz��t�+�hM�!U�zX:C-U��(H����/�:M�c�r��V1����H�95l��v�J5,}�ċ�8���ԈH` P��5j�b��x쳟��r���I�z��+���}G>��O��\���S�h�i$~��;�;�H5*�s`^�=*��K.\D��s̉G]��2DϺ;v����:#��� wT�L�-�TO13]#��yH�f��Cr��>���dI�̙��=[����R��K����A�1���d��,��	N��!���<R�uv2�N��n�{"Q�68����du�U5��8T�"�����>*��Co$�^t{*�vq�����\K_K#60�}�gIB'�
��}{�x�y=x�$jt s�uz��yY]^f�[�����?��T�^}�W3��G�����4�6��_W����s]|�G���ٶ���i@ق���`���wA���#���S�=._�����_Y�|�-?�ģ����O��cG��҆��_>�����^6f<K?p�˸F���\��*'O終��H�p�x-G.�t���rXY)PS�O܇��)ut P3�����hU�S�j��3p��`֣~����W҆yW�u�e�o��L���f�A�:���s,����<��;�s%��������m�R��AB��'�c����;�
�i��V����zZTԃa��{S�O��KI�7X� ?�����:P���^!kɌY��ΐ2���1+	�B9�u8*�x5T��fy[�?C��1u�����3M�7��Qǁ��(��Y8v��1��JRκ\[�s�(����
������Tyۍqӡqrn��A�s�v�
W�n�tJ]�e`�%/��$S���0�=յ���x�7����0E���9�;�Sb�#���A�zcֆ�@1���$5x���#j��F#�;��)D=�t���͒�4v˄)�r�ƭZ�W���>��±�A���~�����#��F��n�!?����:���TN��c[ŽH5NG;eT�M��X^|�E���@����Fj����ZX���T��>�Suh�f;r��Y\�,��C�����zx����0B:3�{���u�pD���P����|�?(������C�Q���K�'�y֌A��;�qFT��=z�:t��pH������{<��r��"���UN�:��|�m��UM��f����O*�����+g��d�}�������!
��-�dBO>"�aZ�Z�w��G�Ş��cG���0G�>tP֗�ʖ~o��g��u������0V6�}�gq���A4x��?w�'���|�+_a�L��.�����xu�Ѓ?�
��К��C�Oc�x_�OM�����<����?���Vf[����n�u_�sn�M�Y#5�h#E���Zd&�v�]�{O�á4D#��~;�Ya���l���V�x��<��F��^�\d��'�sXɩ�8�%chrl���>��N�>��ݒQ��>�z^�f T�/}��T���G��G�Q�Y�+��P>�_�7��/�{�ͫ����l,��� )��mo�3�{�s`�{8��}p!�UG�!�A�_O�"\�ti<� ������{�$�VQ1�����X_��7���F�a��(aia��^��q�ك� �u�ג��a^|9��5��j��k�d��=��Q��R�vPVa����5�M(�{��)��[��l�TQ|`=^��!5�ϸm�&ൡ0R��dY�ѳ�g�#�~+�p�2~R�Ha�V�Q���7�dR5p%��!��rw���
�A'���n֚���������7���)3�D�@��T�=���}�uE�&�|J��i�E�$<zJ@!���jN�8���&��"�W��j�q��^<X��;I9	�⨩�t�}�5��D8� �X�҄y1�O2�GL��1�C�C��^zLP�7��#*=t�lo�0���H�ߒ
Qn�jxn�f����$ǥ��c[2QҐ�a��!etC��@�bKҼ���C6ey#��Mk����nn�X7����M���9�� �����Z���g��٣���P3^$��s߷8�Q�
=�`��ĳ�'��]S#rk���^�ꐬ��Wϙ�R�47Yϼ=�^�O?�4ے@DC�T�V�7���Sr��Q�LU�j��Z�/�#��E�����W_�3o��1��N>R�A0&����sG����^h��ӧ_ui�8Q��gS��;JU$������AHÇ"֧c)�r"�p?��w�;�|T6������+/q���.4b9��<��wɵ�5��Q'�XN���p ��Ɂ�{�Ƹ�Fl�~�k�fܗA�:�(������{]����7�E��G�Y���d��\�|�j{r���SG��߿pZ��)���5)�$-Z��J$��=p�$��` �@�k+��N�U8��GY���GA�[5�����-N9ĸ4�뉵e�ALD��rggKΞ=+_�ҿg��#�~��0���ݒ�ޓ\?j���}�ϙ�}�Z��A@�fC�K����>���w����UD������hT��jy��{�����~�,�χ��a��쇭��kC^H���^)��ӷ�[y�Ջ<��(�]�Y����3���63<���e�͕w�����m�����V�ӓ*�h�+���-�o$��ߟ��e�^��ĉ�(	�-�#�;C��%�-0z0\0�a��1��i.�8E��0x8���FTq@r���7hY��~�1�;��+�H�_�铱y�=߇ �JƏ�Z�8Ti�#�����qG�|H���-�j/TC�i`?���P_C4��3^���s�!�����=�p�b�F�ߙ�u���e�;�B��~u|M��РW���i��^��5���Pf�[��oI\F�҈}V��k��9�>�~�Z�E��ܷo�3P�� �]iF��胬C��F�VúK"�q����&�C�����{�q���	���Jr�����mطwQ��ߐ5��!��/�8�ԔLi(�m�ݤ�G�66�w�e�F��5�>s�{ʉ�ψς60dk��@�� ����:3z���@�"���b|)��;}Yػo��k�c`�A�G�X�0�xMe��AaN�ዯ�,_��5��f���G�O<�qy�>��L�CZw��]2��J?~���۳����~`l	�̰+yĵ�Y���	��j�ȸoP���ؤ#	�����$�s��5��j�/�������$��3��{���Q��F�'x�����Jv���z#9�g����|����o_x~|�+�
Z�龱�I�k�Fl�þD�����k�<0б��7��n�	��oi�8��t2R�С>��$Ѫ�ױ���F=���+_0E��֔~����F��3a5�+3s��<q����J�pW`�N�c�8�J�g�P���#��ɯ�L&g�c\�.xD�$Ρe�pd��5N�,�/I���h �G&-���mn�[��M�L}-YT���a���i�F���P��ʅs�E4��z8r�Ӑ.u�����i5'T��ӓ�����+����S����A١PÏ��6z�us��FtE�G ��$MEl��롎����Z�>F��ܥ��
Y��'�MW.e���]gܕ7Ν�\D�Ha����B��3� ���"����KׯQ��$�&�͍-��]G���Ы��N�܂������8����[��yW'd^�׫�*b�~�r*�{��s���C��,����Nvص�@��L����Q�N{�d�c-����s�!'����z�� c�5��?Ĕ�	��=L�&����N�0� Y����lv�r��%I�ޯ��Иu�p2fi|@$������^�L��7�q��v��yy�嗤A��T�j<�cUc��=��N�Lk]]�gt����€_�(sqN(ҽ�N�i:=y��$��X[�Κ�Jl8�,�9u���GI���~�-Y?����?H�R�밥��Xc�`sk}|���6���4emQ��}���aG:1����!ǻ�Þ�!����$p�� ��2�.G�Z�8_�-��ܕ�Y�T�/z��,օ˸�n F��Ra�i��L�q��1�3��DWu*H?u���>�KD�|8��1�8��)t�֦kQnfq�$3�wf��`0h�P�
�vl�D/�(&�6M���>�Qo��޸�R`HA�zT���*�ᡅo��u��K�O�}��Y������E�D%�F��to0j6k���F^����2�l1L%s�Z�" :����6�9��G(�U�����]=��t��u������}ț3�l;B�^�a61�~�W��R�v�œF��4�to0t�%=x�hʇ�R8љ����)�o��y��㒡��шi��0[�h��P�F�ͦ���eva�m=0pb0D�baȌEED�"e��i���*r��oO��qw���-Fx��������~{�}2 ��x������k��w���e��F���l++K�`��������aFY����/q]����߽r��NݺC�裏��0�n� �ŇNvqq�Y\���}�+�寻~�;*2�9q�&PCk\�d��vd8p�8g��Þ�ٳg��p��w:�P"�@�@��ߐtK�0�@7VǱ�(}��аT:v�ˊ$��O���\��kZ#��U�n��c���C?2kz�о	u�7ϝ%����;c���{�=�{��VԵABľ��[�/��q^��#r���c���������k'hC���4�H��5R^�{{]�'HS�u9��<�?�kvFL����u��ž+Í`�=�]9 %�N�F�9>�H4��@q��,�`MI��?(kb��0�~��� ,@�@-P7J����E9����P&�(t���,ߐ�z�3��z�ظ��kU��5��-''����wqD��a0ĥ��N!���;e�%�{k�!>�Q�h�I)A$����u�b����X�ؤq����{���88^y��]Eo����o~�Q�oj$���_|��?s���tC�������y��ב�GY3쫱�p����g�i��ɼ�{B���=�ً2�J������K[��o}�;�G�ǌ^��IK#��o^��ո^�s�P����6{ҟ�������?�ȉ'd}uM���g���kd�c�4[3�c�q��/�Փb2�{2r�d��c�:�$a�v����=P������.�s�2�h�˫�n�5��!|Ҩ{��W_?�,	�dkvN|�����_�Y�p���-�5��(�D&��OPC�7��͋�<<�u�SÁ��b������%K�jP���QC�xԝ��s��d��wت�Q������H�=�{�[ߐ����z7K6
��wL_��*��A�����j�j�a�������K2#[䤒��B�?�u� t_�:u=�����l�h8@|G�ߑF��kk���*}��{�G��NV�nU��/�㑭j`v�g��F6�{��s����J�Y��0��욦��4�����������dt:�zF�0�N�m��h#�}��]:~T𮰊�����R�hܲ�Q�`�����2��&=�^���GԘe���gYDm��]�]��;D��=�2/r���Bi�pa�^0R�1�4������lkVz�AIԨB��(Z�n�\�kחeUE�A�đ�\�Dx�zA���0����`����{�uh���k����3����Q�� ��s\k�;d}uI�0�Ψ�#�������>��9�@�>�w�~W� ��x���"�m���������)[z�]�~����j��=,	6��t�slv7�s̛3��V��IQ��E�}��A��:%����W����1�"���tո@��̑����ḾrA��/g�3\V��;D|[�����C��t+�?)C;a�q�59������/�8���Ϊ��L�O�*��T���<x!l��I��sQ�2�=Ij}���H
���ա�^9"^���_�+W�;e8��"��5``��UN#?��W._�����F�!O��{Y�Y�{� �d�S��=�Iy����?��_�.��:s�>�i����y��S�T�DC:�1�G>���O���`���'�v����CH��C�0��:���՛j�չ�E(	�� @�[8��O�9f���w�s�K�$Ȇ�N��.�fe��5��Q9���L�FK#xL���U�����!�Rj��4*���~G���fZ܃��`�a�'bO��N"ǫ�Y@�F��:��}�S����H���:ǎ�Öέ�5
���b}#�`0ZђI�h�h[�7r4:BG��8g��8�A�@��̱��Z���N �sA��d�w��E�]�$�]��;D��"j��� -k��Hg�>�5b5� �%��9�k~��1y��#�ة#��W���`:�����{��&�^����hĎZ#Z=�ȩ0A�+��2�υҞ<~�91���'G����T�B(�ax��$-������#�~�U���z ���ғ�A��fcc�ξ��ߒ%|��B�;�X�#W�F�="&���pS��;%��[�k}�i��v��K_�Ӷ4+z�l����믱�٪˦��gސ���K{f��KKK�A����	<|�"���o�ީץ'��qS�mO���g/I����=�:뛮7�:=�wz����	�#��m^Ǎ�E�$r�� ȉg�;�6B��}_�ԅN�u�Jʴ2�<|�z�<��<َV��Cq�f���P����U5y��$K��� {0�&�q���R#�HEJ���Ww�z�4��g��zW���x���=���6���Ȳ�pF�H����l9`��BlF�[cC2����Ad�k���E�uk��ѽ �G� J�R=�1q���?%��`��	����$��Q~A�����NG�����.HT�O*�V;8P&t��~'�3 q4�wd�qA� ���#2���u��ޛ+���Gn��˪��	V9��::+p���FD^D9?3̈���߭��
)D�s�����Q'#?�Td�"�*�) ����!u�ɗ�n�իW��}�{EǑ]�<��P��.��\�:��>�2�x/�>��sY��I3��nG�mJ�������ZR�<��3�w�b�T�b;wĔ6�k�J)5�^�9$��<r`Q�5+�7���� ���׬I��1�;ۑ�3��{j�-��t4�F+WH���+�yQ�I�����Fڨ�Av���~�=s�	!W�᠇��ֶ|��`mmH���mﮭ�VH���x�}��pz����w�یv�T`j��?&�4�1afNC�"�s�='/����������)y_ʍR6ַH�9��=�j�&E{Q��p�~��'�Sv���w�S��թF+��z�`[�2����8U�j^#�g�� 8/q�C��P?#,�tA2u�7��Q���aM�C����U�)�Q9���P������vv�����h��O��H��wȦ�'�MͶ�ة�Aw �1�^(O�Q*)�� 6���RgP0lM���A�n:�����p�￠�����&�dEv�e6���2"4�}���O^{󒮧�mVp2]�g�H�z}gt��t��uC��5ɫČ�j�#]3�Ĕ�m����|�;1��.[��F���ְ�����Kv}�a�s��Ύ�q#=��I��#��5Or��5}��e�`d,J#�ֈ�-7���t8ޯ���˫���w��Gz-�92M�:��'	��	K/z���Ϝ�Ca
�ͨ;гh��ٺ�}ymU^x�=_f�aPs��wr���x����� v�QG�z��Qϡ�R�����p�V�*2����ڳ�
��8s���{wG�<΂�Tɒ��N&
�%�k�n*�pW`��A�L=��s������}A<���:)O�<&jೕ�ԍx)fT�I�	�0E�N]8vP�m֋���k�������0�7X�Yz��0�a�cV#*(iޕa�iZ���u�-b�
R�dAO;f)��Mo�=p�Ao�d]L5�7�V��иohT�6Dh���G6��@����yh"rb�0�z�crՑ����pߞ�L��tf)��	lr8T���{F�z���V��ǟ�Y�lj��H�M
V-�gB����`��K�+D2F�j�ȉb�\ ���:$#����H!��:b�-�a�~�mw��8��x�U�Z�;�up��ǽ�zt9Xd4�E�zo׫~�Vt��6�꿷��;)����EDYw*X�����a�ú:��� L�]�bX���![�ϭ��l�:�j�4P>��+R�h����̴� ?�?ec��AD�%�ub>mh�זdk��#˃:o���>�\d�/����l�r\��s&��!^W�U�﻽��n
���U#��;sFZ�n�=�߽�Q�~�2�3��Y����`AͮQ��HO��U�V"���<d��@nC��'tڑ�@���9��"��y���*tB�ƕ�
�<�=�s<P&��Z�h�nӏ�s ����:�_��7/\���_��wa^R��phqw�r�u	�'�gE��=�_\`K.�3�W�Nq���?���[�؇�=��+z]z��D9b�K�FMc�8�À3��>wvI����
N2qLO�=�`��}��ay��c2h��QGM��l�a����a8t�QO��{��%������E}�kNPEC[W�e98��L ғdO�,���P�E�|��9�_���Y�8��g�k�[�GT�9�	/��3,b��a�PWg����K���~G�߸�zgw�/��u��Y
F�8u����~D���1�`�Wu�s$��ϐ�D[�vh�!+���Z�c�X�ыN�JvA��eh(��MG�����y�!S�y6d$8?ߡ���>��d�i��t���"%6�Qa�6ĊY�;n���E��J����\'��I�]��O2�+�ާ�v?��S�7ts�>8
�Q��U���w!
:�x,c�]߷��]o��T0�[D�y�K�c�5*��H>��C\'����F�� �w]���}������j'O���WoJA"]{ssNZ�pm�N4������]�*�k�c2V(]]�tU-����U�bV� �ԡ�P�~s ��}A��A�N�~p@�KH�B[�>7��Q�h`̏ѐ��A�� �]ѽ�	j(̈́3T�Þ�z�z����y�49�h)Cڝ2��"�j��k��օ����"(���'�:+�f\��*z���w^|�Yt�D�+ѱ� �V��/�Ѷ��o��2�U���^L�"(+�r?�]>�H��V����>/�i�Ӓer����%����^d^���e�A�Cd��ǉ������%h��C���=�'��-�ΙWe��&��e���Yzӳ�b��}�0#���uY�ؔH7����>.g�_��`�3U��:s.	��Hq7z���%�_G?/�0)�����g;q��s�0�+Z��=t�='@+�Z"��%��\oo�Hz�q�!��ڊ�jy�k_�uZ�9�z	9`�^�tQ~򧟑������/�6W���-+PYC�T7���0gІ�%�w�5�A-�N���z_#���S}D��Z���7І��V"��-�"���o�#C/ЪTs�R��H�툽�ҹj�:�:���?��A��H,@:���ގ�]E/0dN.s�0|;L��� �Uq�"U5���wfR'yGc�9�C����[�Z 
�z�u�#r"p]�5��\T����=m7k\#�J��������[Ő��udj��g�,����^�ɹ���-�7\ȉ��H���\��Nb�b@<�r\�� �j��4�k�=�E:���\�|I>���F�����Ѝ�����3�P9E�6At�CYv�
�^t�P���r����L�?��F��^�h���N����#r��uY[Ybv��a,}$�)��k,��su0�&��u{9���t�v��������A06���\'�Z\n��S(p%38:��a�Ɩ8��� �1���1qkl���0Q� �RҞ+A@(L�4ģbw͎:������b$�PT�N���׮�Ɂ4r�8�����$D��n��"�c
3�e�N���n�����G��JjT�$__V�&/<�H#� ��{�*��D���>�<��G��/�_[�a �ZN�)\��z�,z��5��7�7ds�s�Z��d�z��us6����9�E�n|�G �n�����٬;��8�p ো�n�u�XD���=�a�}��-[0P��(���E��H�}�V��59j��4
���jW��djl�q��mA$��W/˪�.Qp�a��wZ��[[��smGJ�/vx�"��zІ������]�ѱ�	x��󲡑Z
�r�5y�<�n�i��3������>���W�G�/���V�;�+5��>_D��o�3���Mt�z���k]�O>�8�X�C�B�:,`>�[�硍V1(��SN�� ��?H��)�/�*�{s~�F�=5�[�����T؆�1!DC,��w�A�q�����q�[Ҥ9���;Ͽ&AIؘ&�C�u�b�ۇ?�A��?�3y��e�S�{��Hs�#�8���mb�V�de}M�<��n����r]����3��4,:0�9��j�c�u������1��N���1����oʂ:����Hרm�}Е3J�őe�С�E�nܯ���L��wT6���UR�3��#�r�_�Ǟb�=Dw��a�"U��s��9y�F�|^��u��qq��k
�(M�c%��B?���a˜����!���a�h��4��+a�T�W�"��3�w����iR�B�ؚ8�q�&ڏ�����7�1ZM��}�A�y�� I�!@9��9Ҟ�deYV���a^�< g�a�c�M�9�~�36t��WyՏŭ}�3����Ƌ�j�А�{�R�N7��@�#'�
�Ԧ��ƈ�?`-���56,����_��~��g��ߞ~M�!����I��ξ��5��Fl���.��]f�;�Qw��Hw#�ό��<_���;���=�)Q��r��]K�^[m9s�M���!��k�CJN�:P�N�w>��~�}r`aQ���O�=����R6����!������)%�֟�SGj���e��!�F숇h����5\����%-����>�JF��������%���V���魃\*��� K�^�A�@�ҟ��^�Q&��x����?$���'�Ƈn�y���Ɏt=����0�����J�92 �{e�&���*]���-f	��dpp����j����+�Pc�AE��b8�&�a<j�icC����勗��O >wp�>����Y����K���<x�qy����ڥ7(����������F�%�!�ip4@��N�����6+;=��@"�"�Y�+U��I�.��t�&�w�P��qm�tͺ}
��T�������3F� ���-�kJ�e�9�ا�YS��"F{��9c9޷�E�����ɘ�:d��_*���s
Í��yud�r�)Ҁ�]��Y��ުI�y09ʳ�����~~C��!�B�G:͂��"g�]�2"˗F���0�~�`2*��.����V5��ںyPGG�r�Y��=bF��^it:�a�
��YW�,�p`�|���H!�p��;Sk���`�8���ƌ�t!���Fn�@�mJ�挼q��l���8K�/�t`I����)dq��x+��ǌHB�9����"3 Ͽ�:u<ݐ�(I�ÿ�ԿA� ���i������WjDA<c*��]FĐ�:,Z�P�w��� ��	?z�/�k�b���M���)��{"���k:�᠏���"x�;d{F
5r�s����W?/�j\9"����\�S�-�?�{�o^�*{��k��_h��%}�U��epKD��H� �6�Uy���2��8����C�t�o�-�d�O������]J/���V"�����נ��L���;%�����ӈ�3����O��������C'�ˉ#�d����_����n�HA�����)(}�G�������d�J"��ۖ�K���N�=��9��_d�%l��^���ih5`�����s�����	��?��<r�	����C��񁯍o�Y����-�(��h�z�+�����Ak=�a<�ǡ�Т���?x��os�!�q�T\t]�9;EQj�� כ�T=��+�]r>��;��̂ĺ'6u��MZ����~u�߸�½ 2j�$<�O�k��.�� r��Fz¡
_7Gʜ��DO��w���H" Jd;��mr!J��]&���3�Y:���#sa�[W��B����T��:����]5���#Q��)e���s?0�,�87�|����]��;Dؠ\�36����8�6"#:�@;���7טΛQ���i[��꡺t�<��,�~�FksԥU��)d�AO9�<Wc�f�h]#J�D$�#�4ݔz\'ZK%����Jz��m�j/
���t$֯���'1�a/����!)�̑������>Hf���CϮFTHy��H��*�FD$������/�ka� )<���jC=Q�~�j7:d�����Ѐ�VD-�hꭺ���!t hg�b��^���ɟ���ސ����c����Uչ�E����!��y�	��'������,SҨ��>�콼S�&�������M��?}ӵ�X�K��Aq�U�iu��?���w�sD��>J��N�";�1�SdA��ݔ��O�<�a)�������yM^�{O��g�y����'z-A�D_伣Ǐ�aΑ���t�7e��Ȧ~���˜~7�Q�G�����ҫ���*�W�7b�{1� s4��˫����-y��I�T�������ɾ�^Fyj����d��l�������hp� Π��h� qL_Y�P�?��]}߭������[Aӏ~�=z�4�ݻG�f����)Јy�����'g�?��G�[������ݑE]�I�-˗�K<ۖd͇t,�}����s~���o.�z��E�~�:u.�XS���\�C;X�7��H�C���A�Lf��A��z5]�]e�,���^Uз��%��9'�˳Ξ�wE
��h������S�ck�&��y8﷜�O��	��#Ix~���Ĳ����#�n�:��$@��%-D�h�dV1�yI���Xb� �/c]��ٻ2a̰3�w���e�*��y(;�o��(�C63j̇��\t�b�zזo��B[�!	l�x�5
�f��Lp���$;#N4���t�3F|~�J���#�"�yD��\k78�aM�,F���P��V�nT�9t�Y�Y8J7*�Ќ>'Z�
��S��g�x�ԟ�	�*}��$oUƫ.1z���Y5.=&<��3,�a��}� Y�%�-t1"�p<��V��	*v(� ���ܑ�;�p0���#�Z��pLm�	fa�0���;���T>����3)2Dò+��{�Nd���X��u_5HY#]{��)9��s���%�IF����c]���QC���~�M��r���шx��5�:���xN6ז$��9��P*�nI9B�vS��^~G��F�1��}MN�����M5�_���~>�Z��J���8�(�N9t��8������- ��V���r>Q��[�\�������\�|�S����g��'�̿����^a{!#Zj�ǼL�S�;/�BÄ!(H���
3�r��8r.g�iQ�ߩ'e����k������x.��R��F~J������="�h��� �.�lГ�M�J�Gl���z��x�{��O���:�.���J�^8�hh���D|��a,b5��;���������Dk���r7C N��Y�q����,&j"Ǘ�p�i�$n�a=��.��,w=�� �+B�_��&	9+�kH�Ȝ6{]�̓���&��Ʈ5#�"�i�җ�ސ2�qsV�6z����ڲJ?m���^���xӺ�t^�(t� �����1`��懭R�{�P�C�����K:� hEA��t�ņ����.��H�ii��#�xcVI>�ΝDd�Y\�6{Yϴ7~�[��|84�<Eξx�6�H��j�o�d�"�s�_�=�F;��~+$v�42<zbkܪ�7k��!sPi�$���h�Bt�N'������}$���(uS�HZrƁ_���e�t@���u�
�t����X��/�1(�����P��ď�t���b�N�,�/��n��f��6���ՠ�demE6:�����D�>�`��o�m3]��`}e��aH)�<r�r��%�gѾ	#؀�HP��B�a�ݝ>u2
2�"����$Y�������B���B��dWD$g.^���7���y����ǩ�w�����РC���$/�������r��Sp�0n��{�������Ò�o_���둼y�<�5Ў���a�1�~u��{XnO���R�j�������S�o�3'{�vh%K|� s���р�Kٰ~.�?W�b\��@���o�2ލ�Yk����U�h�ϼ
�Dۜx�]�c���:1��w���Q��
�����{#
':6�_"�USw��p��P�A�� $OA]XDW8Ȯ������1�-��i�|�)czp��3�Ӓ���\"�)�7�ܐ��c�^���>/�仼�5X�09�%r56����������/8b�	̈́��*~C���YHu�Y�D8D74���ٯ��4�DJWdS���Oq���o��k����S�Н������A���7��*h NԼ+��ȷ	!r�v�����|�9yף�K�ݗ��:������`��+���8`a� i���#�����5�o`�H>�}r�*�ل���JŚ<���G��.D�a1��~��:)}���������^M�z�*'�!�;��ޘa����ʊ���iٿ� ��q�@���"�i[EK��]5�+r��5f�
O�;~�<z�$y,�}�yy��F�x}�������܌�<q�|��ǶXc�q��'!:R[���_ҩj�!�K�BVyZ�[�F��#���I����B�����l?k�+o�!����&K���{���ި=����_�:-����a��f�� ��P[F�����/I����Bvz)ʽ�
�&J�^�����'�S9v� 籧z͒��;�\��Xa�����X�x#xW�v�����V/�c������߈�J|�v@ ��9��ve�%q=�Ϡ���rc�sߒZ��A�5z��>��4�X�&tg�w�YO��sDn�����I�}_z�U���)Y=�A��0�~�����I)���yY@mb��/^�'�I#n�pԕP7��'��^����"��hpym]g(�l�޼,Ͻ|Z��4�D��
=v���&f^<C;�	5� r�rH��ob"@��؊ҷ�UQt�;���Y��&txd�N/�2�i����셯S��ܡ2��ǌ�}L�xWT��O�����L�m��a>����p�'�v�~�WC���O�������K��a/yK���NWR���s����Y�}R�����H����='���3�Ѓ����&��/���;�Ņ�[È�kutF	�B��=ʈQ%FoctFM���(��D�aQ��}��ι{/��~�j������W(j6l{�y�ъ�摭yb��'o���9�^�Fj>/�N����?۹����;e�)X��7���|�"6i������I�����֠{{�q&o�2�Z�9`�.�f��
�B�+�U��F{:�Ű�L�-2H~Eu���O*�TM�ͤ�u�q$�C�ۢ�̠u&˟�͠(�������'�[4Ny���mX��o6P<Z�$)xݰ8[Ҧ��%i_�5�
=��f��>��J�p���쉚{Π�N�nkK���j7��_�u��s����X�)1=��aC(^"�8�$��ot�u^��5�`�=64}��2P�R4�����~�հ؞0�O���2I�P���Hz�T��H�$S�lwB�!��6�_�0!��������]�۬��{��L9�̭��?^�{�nN�����v2-���C�E'������_K����6	�'ᝁ�������W���T�U)o�-g�ɀ�R͡:�B���{v^�Q,�KY��w���,�W�P�w��<ϒ�+GaW�uh�e�3�[Jzf�q���rM%�	Z�{�N?#��!Q�G�egE����v���̪�E�娢] ��/7]=�'�W�k6���z"z5���H��������q���X�l�� _���}�;*b+&�Nj.�pb�w:����������r���p񴧩��LA'���*�h��j�0���p�"�����}pP4�M �z*�y��%������m���S��,')\�9��@�e�l�=;���#:�k������w�^�-��;���[����R�o���G	���p�?�=�,{��T�А��왵H��Y���cWFRul��j�y��%%^�SEyL6AW	�o������m-rx�E���%�X@���y����o\D��L�-ZFҤ}�Y��y�?����d��;��(�P�u���l�����LV^���	BM.�C���6��o
*��1/b�D��Jߋǂ[���e�AU����M&"�O�_�qeE��_��X�]=Ȼx)ͽ
3#���[��"Dݤ<̎���΃��'X��ؑ�2h����n���x�u��0����h��s�(i��]��<�@Blh�,��N��p�� o�q\M�6م�l=��kai�PbY�?��"e`AR�.x�hW��L�;�+��NrN�� ����ʲ�	Z���rb������@�L�#��i����5~��$tP{��r��h|e�&�ōW*������v\��z!�Y�ͧ?ݯ�=~������?��S�m-�zGDnM��`C�x��X�񁯏�u��,��u��-�T���<z���L����2{y^ `?hB��Ey�sm��+KJN�=����*�LUH�a�PmX<1=��.~�($�^���I�Co>>��TX<����y�I0t� b
] &�O��o2��iZ�Q�����3;����˰�(���C<�1�i��w�
%�}耺���X#l���Qo#�O@7U�4��u���R+E�	,��rSFQl:���Wz;�j���j��N���7ݹCu��3'��'Uk�a�X]�$e�I+4�H����f����`)I�-��n�}ZEB�N���oG��=o�����nk��KBR�pY'��#���Cgo�j*�?�)3�x�.ʙ#�r�Xf����(z�P1��cw�����R0V��E]��~Hٯ��g\T+.�s��� d�⻜�)v���r��9���ώH)���I�k?؊���g�.�3�9�\��>�g��۝����V�y�>����}p�]˹��,�nC��Cg��`�\Ӆ�Ĩvؚav!�ɯOJ2�/7^���׹w~/�Z�� �Z-�Pڗ)OE7��z䶜Q�� �2���O���z�Y�K�~��G�&[��b$���_���:2�����G�N\�P�f�y�&]41��Gԫ�M�WZ�R���\����Gѱ�a��2����gp��/��$�Juҗ4BU)tz���e}rg�F镱�>�~��V_ܪ� ��؆MP��;E���V|�0�׍WQ����`9\k�Sجe�.�9�~~V8��,WM��d�o����t���l�dI�_'D��xҸ	�64V��d$��>�7�U��l�+�O��>��<9y�*��E8zq��b�+qR��I�x$3l��r��jF���qJjX���c�$�r}Ԛx��b���3c�u`M�	��� X$`�+�����6����{��`�b��	[](X�܈�n2��<�ý�@ �MF�B�����IB��Sݬ
E,b��g}���� �9>�g6��L�ڡW��ϙ2�`#�.o_n��:xQ֭*��(e$Ga蘫�oG�ڤ��$�`-�	�>k��+����*?ߖ�������f��T�d
�y/�.˼�����4j�A����;
���y�dϵw0Z8��y��������#w��AOݿ�h�e�$�@���؀��������?�5=�+٧TA>,��%����oW���i�O=�o����2(���e����]EF12=��7�����X9u �f!sA����r2G��J���r���*����:��A��w}L�ez�2�(if��,9ƭn��� �&,9?�b]�� h�UIOH�8$5�Xz;�d�wC��8
R��t��Y���d�CL��&E#��f*�%ɳ�U����VndЦ�i��8/T�̷8������]ƒK,#z��F����$�������.?�2�f5!̲�7P{�|�*O@NQ�(�.��O]�W�o_�ȇŁ<�d}R�'��Jx�r���w9�\7o��i������y�.�}��լ�
g��9�(�3j�+����Kgpn�������{�`���B��+��e%^��M�J�47O����iR�^r���z����$fH��<������8�S�#�g��=�/�5�d)[1|��,I�*k��<Ѐ�g_g�)��2��8*� 	��p��J���</��>q�-�5_�%��~�e�U8����t��Ҏ-OY��f�9�u��� �S��3�c��?� �	� 	>+(�.�U�����uÿIV�6uQ�ͱ�j;F���iTTg�F���O0�X�9�)�N	��2�K����d�,� R�|�5��/C�n�,�΍� k(�,+�S&2R�D�.��+��aُ�6tۚt�'HB�D�S/�e���p�����t3������g�o^��J����r	'�J�䱎w Y�������L���@V�@͵x��%�j9TAGH�i�a���}HD/�(��)��Y�����/��H~%,jQ,�w*1��8p�=��%v�<���XZ�60�S9lt�C�
�Mxw���f*�s�eK1o�L�3�r{e�`��h�1��|�Oɠ�р��2�#��yZ-P ��QDI~�W�'�UY����~��PM�\�OH������� TYAߪI(	�c���6
՝c4kW�����'�L9�b���k����Ko�xȚ}o�p����Q�|�Ñ!�{�{D� ��k���f�A�Ǝ��Be���%~w<��6�)|զ�Z1�n'���GҴ�_���+x��)�ј�Xg��0�)��b �FzP'G�:s��x�%����l5�͘!�/a.@�O��<�!2E4A�r��H'p��vw��p@�3�#c²d8�C�b_�];�s�f��(��CAA�?�o%|e�dq��:�x <���s۹���K�	��a�RzY����j���.$+T�V4�h��{�3x�XDXi��A��>i��p���{h_� �'j-1 �e�{b#�O�������A$���\W�S��ؕ$c���b%U���{(0u�c���W�^d�A>�VK"L�Z$��u���o���=2�vk��JM��M�A,A��� S<�T�-���:vfya���n�i�j3R��Q\O�7{G g~ӊ5�ߎ��汶���B�]h&nC�j(씼H "j��'6�*�/}ؒ�y�����9`�|��Kyn���*�h��Wӷu�,ej:��U�w7��	2�,�Dg��-x,0w?d,)Z��(۠Cj�J��b"��fԵ�n�+�vWah��YN�����(F)+���5�����������f7k��Țz(g��<B��l�q<Q�d̶d\-���T֦,/�|�QT�z��n���iU���Fcz��œ �WX[!���2C_�Fp^�~���ڣ���b��TD��i �
��׀-�*����s��^ow��P�=+RBԖ�� ���Ȫ�kB4,���/`I��|Q�d�����%ex�_��B��G����T3��q]�����<-H*��ٳ`�т�<}?�"�+]G};���US�S��Gx�T�X
0�7�f��4<��W^`��qL7M���T��-VO�l嘫��g�6fغ�5$B�4���Qa�o\p�4��r#j��ぅ���95�0�=j��ϱ>$��m�r,6�@u4����J��$ }��m��9���\�Gq����\�,���bޙ&�~1�-->��
׺;�s�����b���S%�6s��l�O�!$����m��]3̭�<��ԥ����3G�#��AP��3���U&��,Qm���X������T��iM�~�^c���?��B ��U=������wA�E^�{�:n�d���uP�{֢�0dg,w"�~�O�[�ww�|P���������Ո�P	C"A�(j������=.-�,�К�3~,�$w�(�W�@��2~��5&�s�͒�ò�M¨
��g��������A_��Ϋz
K����"�p�󭖏S͖�13��V/ɠ�7y
7cŀC���56��=����#�Y��U/%��M��#��}p!�m��[;�k�L�9�@7�8g�Q(q0؞�m��<V��7n7�RZ8��vp�'����f9�х�nfh�>+�V[ܧ|�į���0��O�$Q�:�9������g��Ѝt3��3�ۢ&"�?�VO�&���+7�V)��S�"��X?S�v���M�E�Z�e	�=��M`^��|}�u��p{-/
Ϊ���cJzu^%/���{���<.����s��ͫ&�㣔39���B�����(�6�z�g'K����I�L���$&����]�=ͪΐC^x��U�XA�o�s'O������5k
�@���}���۠���ҧd� �N?��@�8}`������Zx��8ZR�tBO�� ��$����G��v)V@�1P0���i^ؠ+�����ږO�xw��6��͛B7*:���7!�<�����
�n�D�+n��:�Z���7t(����wsZߏ�YD�(j{��n��o�Ne�.�I��L��b����Bw�H@��YX���b�Ԓ�](��7�����6XHP��/&* ATh{�^n`g�BFKn!a��N"�S��x�_?���_�]�he�XԯX�t,�F�W����� �,[���0���]OI�O�p�h�S��|Yi��+
���;c�;��Js����M�v����J�_���oPO�i��2(]��h����͸�]��o�/D��6� �Gc�Ld�ݢD#���	{��Z�+����؈>��/�/�/�/�/��
���+����$v���� *Y<2b�
<��{]a��l�v�DY}��o�p<��Jn�=��i��U�ؼ�PK   .��X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   �z�Xk���  ��  /   images/aa6b0e15-4878-4df8-8b7e-ef384cc3161e.png<�s`���>������mc]�ն��mc5׭���Nm[���x����}�H��s�s����U�2  @���P `!�3Dx�'���Z�_H�2:� @b��T*��C"7Im75'K7��7 d�q�s53q�`q�f�}.� ���S��9]z�̷�^^d�ϔ��1�W���쳐��d���)�������<�������X_�~�~u���Z�A�`���<g��6D�cl���?�@d�ݕ/�`\����Q���D��?$��7H?����ԇ��VF��x=���.���=s��K�������C�B /�v ��'����vd`���Zf�#�]�+��%�D9���p��[!�|Ə�AX�Ti}��2�UvG���R�C��)��D�.��P��M#}E�w��TG��l��#����af��b�fo��FR$c�qd$qd�h��Y��!�a��)�/�7*�v�n�0w*�fx>#G?f��� O_����A�Ÿ,cw�3g�#q<��g?컹"'�,!́E���y C8#Y?�~�1#Q;2$�e�2S���H.�$�y�T�＃�2!���j�����ݓ�p���������C�%��b��gL��"m�A�٧t����!��<x��J��w:J%������8)[%J�^fJT������^n¼Ā3���U{���r菮�`�,��w�͖�}���B����_�1�f=���ZORg��Ï���Z_��g	{K�򹗮�%y6ʇ���m���d������+p����=�7�U*Zf����.����vN�I��QN��(;i���S�~���2�c�9��8���MB�g�)�X��8��H__��L�9*PyB�F%��cH��F�m4s��ta�lr-e9�&�_"���u�+�4�zy!�<�E�W�@���)s��}�6�J��*�ߟ��!�߁�\�������Mc:���W�3�%���:��H47Ҁ�r�����"��<Y��u��N�;�t���|���lj��!��R��7�dq���\5W��%��$ R�8�������P�4;g��V�ߌ�"����;�����e=�r�����6�G&/���7a���^�ky�3D{�%E~�"m=Č�� ���;9��+M�1�o$�q���m:�l�_/�Bq��������f��w��Č2��ƞ������.�,���yaR͊��k�`���%��{� d��ۯ@nҤ�ݍ#�b���#M�C~EO�}�\)ȣ� s����qJ���h٤�}p��#��X�O�Bѕ��ô�o��5l<�'�OU���o�o,\�����xXn������oɓ]i�جPX�t��Z��m��>�����mo��EJ�tV������)d`H>V�?��e�������J�F�R�`�Wv�|!�eu� �/�E�����?��'6#��f�=G�A� <�B��{rQǆ�u�S��BP#�H�L=�oz ��W�y"[��/&��/˞��_��nB盥���a�_�P+"l�HJ�||��ԥ��Y��l�s��씝��̐U���>ets(����-��g�s
�����7��fi�Φ>���G������G���7�c����*�jVj/�D�.9W6�h�؁]i?�/�+@h_��8��ؾ�0˅U����ݐ��s(�bZ�e	ښaF�i�S;�,���U���E�J�Z�+�f�Q��fX�A'���83t��:Gg�!�;(�݈��-����G�O7��{�pؓ�q��sp��o�[t��q�-g\5�#@���E��nqg��g��Ϯ�eM'�o���՞(P�ol���r��f�Z�e�Z�W�#/G/v�N>ą�A�<������I&',�-�>�l���<ɋ7�6���4��'{<�Jc'��И�����D�i���y�-���������ǟ O���o���_�7�D>ܟg �Z��H�y�|�7W��+e lw36�J.ح�*T���Y5�?׷,��`��к���O�� ��Ric:^��|�;1�}`�ޓ@�jb#@��<��G"�(��'k�ᖫ9��/ ?xf�41ũ�J��툌D��en�1�2��AvFoG��LnҮ��}඀��PΪU7����QAe�e����J�֧Y�{�\��]�Z��	��Kr���lX�ϡ���G}�����Ӿ�h�?�PF�l��C�]�`Gm�!��=\�G�8������sϥ��h����~�%+�ddlq�$�^M�[Vwa�.�����b��KP�W��y��I��(@19�g�����7�V��������_�k�I�+��f��;/b��}7��o��(8�ѱK�����TQ�ظ�ht��hT����[V���HI����%�5�/1���l?G�i�N� �J`����vXR���o6�=T�W/��T$����u�|�GN�����:7�7ݗ�n�V�n�<�"55[�p��fJ�E߂?y�8C��d��>�:�޵I} H�k�>P�����,;��I9��������7�!<��t���T�B��jk�r!�ա&�,����ս�4�g�~�`4�f.D�
�`�G��\�PN�z1�1S0�||�zœ����h�0JI~�>d���,��m�{v�?tg�n76H~{+k����f���ݭ�0z@q	���P�I��0Xs!��ƳI:{8(�[��
��]�MZ���@�͖i�zE�æ����,�1i(q�@'�0��'CI2�~;��n��g�
ˆ��|��+"�ԍ�®�i�jR��rW3b�?9�+T��t��I��!Lu8N�z��.ض�,ͺh'���L�w��]Q�y Y'L*T�'iΰ���3��l�;陬	�=4u���a?IEb��=��TR~����O���&
AM�"�	��F���}Lnjap8�]��l/. Br����q|�;�`��E�͸�&@�mU����?���]�5�'b��B�h�Ld��s�4���}��"��QZ�L6���=h��kcs���J:X��E�-�u�ku@@�@I�&�0��a��	(��L!Cǿ7�N�fha�Լ��	j�h�HJ�K[���{��!��jl�e���d����<�H������S�G}k��P��ݔ�d��*�1ݷRG�����+A����~_0�|MQ��=�5Ӓ�)�<��3�%~�|���U�_��J>X�H�ݕ6��{�At�������7���@;X�S� �
p��=��ۅ�K��3 j�|s�/~�G��4�\���9�_M&���#-���t��X�z��'��&�wE�����yi�J�h_�aי�^O+M�r9�� �mx��PT��w#�ɖ�o1�k��?���B�� ��S�X@S�GP� ���6v_�΁�!���G#;��n�}�
��q�ޒ_:�D	���&�N���w�@�QK��h��_ϣz�`�O.�S�#D�f�/��
��7P�oU<��b�!�g���㰋Qr����3!��@Y�'(r�Kc�C��`���`����U�.�[��V_͒%$��*�������MZ�dMms�l��i"��=�IE�uby�)�58�x>q��%��.)��g@�s��b/g@1��搤$�a�/�����x�t�v=`j���0	�J��%�\�,z�	�d�[%��1����0���		{�/.���a��|ߛ�{v��s1���]X9~�矝Z��0;#�8n�7{��y�W��Y��o���9�f��Hо�k4���J�Hq�D�֌pE���=�N��F@�OΠD���ݾo�c�5K���v�g�`̲��p#|����,�<�ST�]�ђFJ<ĳCrc㑳h�����1ѿ��燢�=�ӔҔ��cH���tֹ�������w�� R�P����g�m�vp�Z�kV�&�&h�QS/ ���}^��PF�� �8W�Y�.Kȶ�<*����C�����0ԝ�����CL#���1�i�\��P�0��=��� ݧ�m"�ǏڌϪ:����4C�� �y����.J1:C˨������Ԓ��)�(��Q��L>���7��;uy���H�ӗ��V���2b�X�"�ˇm:�Z�d����Ҙl%�!�^�ng�q��@L�^�tB���I��J�U��۫Ne��갴�DH�����4�u2J�@��у�E�.�q>m�JW��~��g<�-#$�H� �)�i��NC2��<��D��أ�8�r
���q�}a��ʚ���� �2K!��i��"��Q�dۻ��@H��"���u�����9 �C��Ɨ�T�f:ڠ|�[y�ƶ��/�#)@����B��1�"c�H$7�nT��9�gӓ0x>h�\�_,`[̴ݗ�w��#�o�c�[\�Rő��e����^m�����+=&JK���Ԥ7bV���a�{�����T���Nh@v���@��PG�Y#O����矢�͌��Z,��]ob�b2�B���!��;��{̵ڠ�-[6t_�2�J�A�;"c��3�":�+��B�ׁ���+� �C�!zߦ�js6_夸����P�l�	v�J���hS��n~emn�I��`�x*�'L{Hvq�H/�^�f�`(�2o,�c�q7_|���76M�="�����:�Ǣ��L�(�wINlMך���^	%�id�i������c�,���j��#a@Mf�{����|+X����q��a~� d�����_}3�m(쁕��[������|���a�P�]��+|q~B������ջ��#����������*r/M�/���U���������IFF��3m��{���# T��Ǟ'�S
�/�z�7�b��ˣ
�������%�	���*5��߅������W-�PF�����,u,�e�8��`�P8���?Iy&dk���6uߚ��_�Id���?Sy�;�EWAR�
m�8��v�Ůp�h�&�N��y���YM�wQ��h.G��BZ�u���YB�B�V�B"r���L{�9�i�%����w�y�@x9�%%#c���>���慺� ߹��N�q�$KB=ʇ��WK�"L�����������7x����膎��g�KPR�a���o�����so�5dcKXu��S��/��U�VNh��_�)��!�}�ɡ��՗sK!�.Dq�;�a�aOc0�w�����Ń�צ��Gb,3�w�,�8����셑��C�Zb������S�2�xn��Z��`Ѐ�L���4���L����"�M&t�C�,�5�5�2��B��Al�
�!�*���B�%��4��o6��O QX��Z�T\%�5^�.w~���MjZ�w�/�����SL3k�3�������Z���.y���y���Q����U��Q�p"&��L|~/BzU�C�wG��Cpk������X-�Uڸq����P,ٴ�S�M�#7E���>�$�ס;���h&���T1�`^)����E'�ӹ��܌�f��̜��Ww��M�U��n�8�i]1Q���@jc�3�
�Z�3�D�ia���kkk��7!�f�[|!��������!r�R����؜m��x���d�1�T��M�8�H�r�s�O�9v�Ԣ���P��	�����"�~�4)�<�މT�������}�RO9	�7�+���6M|˼�wor���u��l�r�jV��v���cS�c�A�T3}�@�i��@~� �i�[��m��
�B�*:|��m'8���XD$�M���V@�z�7�0���_`�� ,Օ�A'������NP*3��@��;�CS9ɕ�K�T��b�P8�>����8Y{�CG�6V=��tk(*��sfS�c��<V��[��&���VH&���ߙ1)��Q��.�u�'Ϡ��Xѱ���5:�K�}m��_ш������ߒ��>_�m���QY>�^����c���)�O���?�'=��p�sT!�D�|���z��t�����!3��~B�C��Lo�If:�Ll[�*"�=��9L�6����k�0uz�F*g!�j��m���0o*5?�H<�ͺ�\���0�3P�6GD���D`�M9%2xH,I�S����qU~w���w�Z�1���(�+x�Qf58w738tq<�� 6c�Ks7lM����^�+��H��~6A����s�gH*�?�X�0���"$���.>5����CT"�+��e�P��B����ڿKj�3�"�<�FcNW�T��dB=3=�50��$�c}^��M�aM��L��@jm��kj?��Ƽ"L�S_��/��1�d��hn�|	���.$�T
��rq���k��vb,���Ŷi�E�x�g���z�U_l�ZT��|M�/�/���nx)�.��LG��B\��Q_�BT~�	J�pW�L�D�r�ߪ�Ժ~�;W/��&=eɤGz�ܮi0����Z��R���r�sR���s>�t�]I[9�/[LK�so���q���F�ʾ@�]?ZX$ݴ]�5@Qo������'���4ƈ���JWt�<b�/t���G��6�����&��}j�TBzڡ(V?}��Ks@�����%�Ա����}]���06�N�XG��$��\��Y23�8Я�'G�����*k@,�nxR��:�4��l�_@�`ޟؼq�|��ƪ���/N\>dYLh��YT���w�9~�ط�x����B�ϛ�q�/i����;M*փ$tˤ�J!����t�a��Bu�w(.R/F��s[�;..��p6�?���*
qq�Y^���?q4�@\�������Q�1K�����86Ig�E�L��V�o�Co�AU;��w�3�~¿aש�3R=�lD�2޹���(]Ol���`̺_���d��,�/�'�R���ɧΞ�WK�
��!kp�ʓ�qST��mq��8<�x�=%M�*� �U ^�Bw���/��郦�w?)�X�##�U�����273'Q6�|v˰�[��&|�;��Èޞ�ٵ�Ym}�a��Ъ$5�;�NV�=��cڜ�bi8|l�6\鏾l
��S����	���;nv��s�?�c��� �9'�]�3b�tL�]�F�zP	z��2�?�>��z��w#g��MprtB�ƾqi�߄����G��B[ 1'f2��;�9��d�y�f�2Χ �p_��T��Z��p�|ش�S���z=θ�"�����"�PC ��$�� �V����Y�������Fp܈NE�۾pW3��R�t���
�]#��N�;,��_������s�+5�[���z��Msy+,�M��21Gĕ�͐����"��j3����:�ɧ�;�ڌ�8q^�B�Η�Yʂ�v�w���Y�e}Bj���v={vo:���(I�69((��/��
��eavAv��k�����S�8w?B?����u��(뭦㏓�	*.^V=�U�u��̐�׿�2�^�5'l�
��:��h�o6������R��ǎ6��il�[�hϋ`so��&��K܅Y��������]<w�Up���g�-�-ސD�QbG���iu��Ȗ��� �0���&���\ $�S	o��;(������V��gA� 1��s�fn;Ĩ�?,�A�G�M�c&�8Q�u�Au��G�0?@�����/�V �'�೗N�!�7U���h16�:�\�2�%q�j��^�Mi'� S��t:��=�{�?�S	�=�u.&�t>#��`�@�z��cP5ٕ��M�O��990ݽ�v���Lph)Df�b���
2e}/�+�O	?ؙm'�V��8��6?�4�5������w��˚Oh�QW��Z��^���ӛa8Rr$�R*��qy��;)�x� ��:o��Vqa4��7� �����|N�l�wxjQ>�N;xI(�������(�H��,����Ư��^��'�ɳ��2?J���VL/��Jt��3Km\J�l�Xr��l����X�������z[�����*7nsv.7�K-d�)�r��i�+/3UJ�>D��l�a)�`�iըRz�*�Sv1r�ٲ��<�"4��a�0��xr /�����v�f���Rk̔t&a��/�-��K��h��5�a�>R�Ϗ������l1s��v���0�xuoNB�w�~�۷��t4&0E>�F�}Z��'�#.T�q��d��'pW��T��W�͚���AMt�|^:8́;J%�-z��
!Ƒ�]���-�d�>���#��c�* �����%lE� �1�]<�PVQ��Z����|�m���{_��(H������t�Z�D�x�VZ��}3��?��%���DB~`�	䞼�/%P��&�M��R(����i2�ʡn��⥋�u_Atl3�W6�(�8�u0��b�<�xb��b	�A]���/�_g�B��m�^�r�~����}U��7rj3����2)V&D����(��UbQ�e�Bf�� ���0ٻ_ғ������7f�m�Y��)�V�$�8"هV��ի�������[����U�/�5�0�@ɯ�~���8ɹ$N<LV¡P[?��n�$����v}G�
��NY�����Kr�2�h�� �A~�c���JE-U��}��{�Yq�6�aƩVR�}��_���H��x]f/to���"�i��m5��$�����*	��@�04�Z�j^L,k@�f�QӖ`gT�b�Z	�^��)MHz
}�a_��o��=|Tb '_%L&���С��b���S�r�6�^����`��@g���
;-��z7iR�<ڞc����.Klp"�|���p������8x7k��*٪���_ǔD?q�x.jn��[O�eܐ\��``l���s겳��ψ����Ud�m�B��^��]��}b�d��;*�X��b�ЙA` NVG��ѿ�'9�;�_1��XH:�dR�Z��sⱠ�8��:��p�->���r7/^C�R�����;6��3rYW���:r�{�%$�d9~��i"�h�]�L�;0=�܁G~	�� �d$���:6V��
�e�����y��#/��0wa����F��%���iJJ�X3G�n��V,�|�v��Y�PWs�[�m��=_�?��>��GFw��ކ����8�{^~��6�x���BD���U�~��[G�N���X�D�N>"���bG>
U�U��P�g��D��[0�Z|9莶�O��1&��V~ݪ8*��L��(��N폦u@����B��DX'!b�B�{_/���_��h G��d��ۚ� �Ҹ+~��M��em����Q|��b<E�}��O&5��o�ZJ��"xKx�T9��Rsxݳ�3�#�BClt�S�?��h��K4NE!�뀯8�=��_�6/~���X}ǒc�e����N�!��
���a������}Y4�Nͥ�g�l�c%-���o�?�S�θ�췵00K�@Nu*!�|��:�����*�UI�;&�By��R�,$Lr1
/���+J��b;�RźD�D�%�N����RԱRi�
����k��sqn��"�Oܷ_~]�%xGs�Q��Z%�B���P��<�{�^����`o�Q�=�^��ZpӁ���
j	F߃L�^bk���R��x�A2�"vU6�Gkpۏ�h��]N�s����
��?�\�}gD�}"ѬqH�%�yl KX&�}f��/|�^��q�S��Ol�^�奉����͠���	+<�~%��N���n2׶vUX&���W0a��ٛֆC0Y�oxF��`T�ƕSb�;�lTLy�����6w?p�v�+3Zv?��Ȼ������'��PjAM�]��M���g�5ˋlL�����:�~��S��<��Ϟ�[��.@a�h/���R'f�7�`绿�A���z�*�w҈Sa+�g���s�G��p�t�������[�+́�=����Y�l�[�.�����d�����hy�i�&Oyg+!$,Y�B:���Q �q'!���J8�Y@�	�ٷN�;	�>��8�&5C��%�`^� ����d�3�祤Uݵ����I�%�U��7��j ����>�``l����\ ��uE1q�
}d�����̈́�E�Y���H���:)n9�����J	N.������3�jB
���ɥGG3��G:��������
%Üq��><�>Z������ٯ�����k�&�M�XN�MN1ݝ<LҠM? ���6ų�!�@?�։=:?�hO�d��@����:͡e�u�����!��R2�"�6��4)�u��ι��.3<	�|L��4��1��y	��ጜzP��9P�؈����O��^i��$qH���=�~p��ۓ�C��B���1e�@	pGa�[?)q�K�C/�Uq�9yAӈ��j�y�՝���x�=%92�/'P���ɳH�H��Z�����M�D� h�
�|�Y�{u[kM��or5[��鋸
����\�4	p���n�w��Ģ[h�X)�Km%��ZU���"v1�d����A!N�HI�<�>�. T;�w����Qq�5�dPg�w0�<�9x�	�~94����;�s۶Jw�_nJY�ơ �;a��6��5xiH��R_� �~.�B1*�]r�E�gVm(,���:�_�D�$hʅ7b�u��q��Ή�m�����櫋d70�]�zmWz�`7��ӦN<D�rvu`�h)ʐ&s!�}]+��0�\I<TJ3ј�R�>G����F�٫��6�Q7�������:h@!잧������?�r�	2W����Վr	��\��:�%��KW>�E��>'���&x5��'�W=��h�v��Dһ�<��W��|~�C�5�3rz�7�T�H���|T��ŝ���9��$.^Y��ˍx[wh'��.K1�;=�]�y���[�+�O97�D@@/� �� ӡ~+����*G���$u�1yf��h��H��p�E',`�䭤�W��1�m��&����%F�-o^8�'���;y�]N�)��-~�Z��5"�^p�bH���(>Ro/���!�\��s����F�8�S�A4�	`+�]7��z��)u\�_��T�x�p����mb0[��������<ȖZ�K�'D)0;4%�P�$�wle�(���\��~Q�<��e�
JɄ�JP�=��p�@�]Di[̛c��}Оq��N"d&%��E,����緉Q8} �=�(��S��_Z����k�_���؇/*�,���⊠���mU%~d��(�pn�l�Zs�8T�s�D������ m�O4	��'�����|A�K;U²O���_�8�8Rrz�P�<c2]����f�T���:�%�FQ���av��3v���{�+lK�S��^����Eu4?��WR�GM�0�'���a��mv��%��vŴ�K,uk/��^^��ߖ������������o�~z��[�g���|{�o����Mt'V���?�������M����F��Ew!�F�Ӑ�y;�X���i`q	׳�7�imD�Q��r��*�I�Q�b�2��ɺ�erd�f�P%���
4W����hʬ���Ho�!{��M#D���R����]�¬�(�U�Zd���Ѣ��?�|]�(Xl�_-�f��2+̮�̧�V$�='�⦹��P��CU�����U�a�4�x�,�M��e�}PU���d���	�O����2����f�^���eW#0��[Xƍ�S/��,g�F�V����orD.�ND狗+�8&3l���3�#T�ad�Iq�~���W����_��p�3������Jz�AG�B�v�������H]����%-�f0-�3mO�+���m3伶�h6��>y>�7#XJ�*w�i(����.��1
�$�߷�2B��LMF���4TƁkHw' T<'+���m��_<x(�JQ�:[u�M{��HdBD�Z?$�lz���`R���o3�ۃ/�.���t.a��'����Ҳ3�H
K�QJ���+�4�)4Lbl#ܼ�ė�K��r���g�
wΪ�T��J��r�β��n�Eu��Ga_���W��#�()B��K�@"���j*�[|�Z�Eg03DȢ:�x8r����T�톽��N��;�zl�x�˚M���&� ��D�݉�J��+&���F�j�6(�-��e�r2�K�Wv���zLw�@��6�a��A�d&�wY��[Z�)�`�M*+��mS�p"�h�K������h���F〱-'o"6�-)	`,}�0�@�QO�#Pr�	t2���rӟ�W�;0vE����%��"�nmԤe�E�s�;��|֬�|�]����S;f}�R�(�{4A8Zq��Ӧ� 8H�rf�x�����]�M�����v|��m��i7���9��ѴXN+dCP�e�JmI2���$�;�p�7�>�+L�� "5�vP��@�"u�X1C��Vm�KwP�9��ک��d	�ʾ(�9�m�E�?PQ�`����r���4n�2��?p�������/�v1����تMo5Q�08�SXy�hXoZ1:���7 �S>+���2��f�+
ˤ��yV\Z�u��Y��.�p�x�PWr'v�G�.E)��v�GGtl�7K�$~B��9	��l�>��h�;j㳁�}R��9$�n{KJ����\����S���2�у���/XucZ�:��狹B�jx�;=�86��<���M��5�ZZ��L���x��,?�Ptf�����tReô�Q�NQ`2S���?�`�Ej�O����Ht;���&�)ߣ�b�#��W�5�OB�euI�}��.@���1�/���8O0As �Td�/�v����wem|*�-���TJr�������:�C8笇��h"j�7������w1�f' D?�{G�xll��|^��\�%{���PO5����y
��TB�l;a>̖����D9��i֗�h~scצ��WV���F��7j&Q�O�d�iE�U_��+-g��xw-n�s���7#1�l����/;�q�$J�X�����T5���Ľ�)�� ��� ~�G��l�;ù��:o6�����@���KF-�^��K�4|��E�	]�3����FŘ|A��id��s��ZNw���⭘�љ�o������8�Ǩ��A��_`�:�B�,M��F�3T/4�������+(���_.&��x|eRUH�O*�2�3�u���Q­���s���#L���`O4�7pW>�D�o&���4ΐ�-<�U�?G3��j�8Y��*�[ͨ�J�����w�:j�6�vƳ�é���6�+����ԟ&R͢W�l�䰓90�e5hlCSU/4CV��#vv~���]6��]%,h�f��]x�Ŷ ��	߅q�\���j΅�nKN�G\�!j}5ϡ�S��oY�t6YG�U;r#�� �<�g���A
�}@<�ߩ.�fR��7ʺ�8|�dùE�o �-[�!I|�WN=C��ݐ0�4�ë����
9┭��u�U%[5�w�/��(\���$���@U'S���s����� ��Ts}\���r�v���].eZ{/����ݮ �a��#���m�[���"����{�S~�bNW�v�>��!����rɖ�Ɔl�5�bx#�����0)^���mw�O}�G$hhC@Bjn�TM��za�<��Å�èk
*f)Z�x7$g�+��$��=N�F�Hǂ� ��9v[u�����U��S�2���u��j]��F�fm��,[��ɣ�2�~^�o�3z!n\yS��Al1ޫ�	�;���3u���%�Y5�~TLgB$���sjA��2S�p<�C����i����֭�[�S��LfVv|lV�47\��挖I�MSx�0G�ӹ��?��W�eġ�˃y�!�OF��6���όx]R���l��i�O���4����D�S�~� N����w.��*{q�݊��14-P��4���u�F�w��]������@ιb�j��@BN�c�Qk��NYQW�qGBB�\����OJK7���@��\u�Sٱ/K���Ȧ�ۥ������N��DD��l�����fj���-!=�¢J�w�Q�|�:c�u�������ƺ�\�3�4<�i�[j0,I~����@��x��˱���Ya(��o�*hu?�39���UЕbn�������:��`8JI0��d*��&���b���c�R��ٸF���b"rp���?���Hҋje䘠�����u�?d��G����U ��L��e�_!k[�6�Z��"��a6^RK��˒��P�g�֝~�4u�}J�����͡�i����1��z3=����������n��$�6���M+C����m�G�JmQbk:�`��E �?a�`�;��E��<}'�@�͓(�2�3��D�|2�)1,�^�P�ǵEeBm��mp����l�����9��4�1M�nè�/��p��,}����~��]���J�����_Z'?�z�ި<���2��r!�F�O5�r��e��_E	� �~�vA��m�:a��&���^��凹kߔ��`�s7O}�����|F]Ҩ|�16+O���H�!`t0�f�8����͇p�ɍ��}7�]�]�����&�vн{�\��V8n�����̍��B$3l"��n����������Ǫ��a����jۿގ���ӫ�˼1�8����%��hC3�ʞ���Ǩ�{�.O����T
�m�.f��	T��]z�Ư�f?��}qs��� �n���:�]��fW��b��u��o�\sn�~�������C�7?���7tP�Ok���E�_w����*S�����6x}��_�:���b���k^W�oN�����!+{`��!�`�=�e��}��7�CAhh��y.�^@����B���:Z��3vS��T���>7a5	i1��r�}��Oթ��D	=*]��{|�q]P��s�'����@^��9�F�~t�xTӚ�� V}F������e�C�����z0).�;`	��_p$����^M�6�|�@jNg�"o�������\�0�>�n��.،_�Qtx:R��N�ּޯj4�� Hu���^���I{���u��^i�Yk��7_C�iE�`m+�8��;>�!Q����,�9�[��o�]���j�!{�
E(�]�\�F�v��#�A,�Z%;�J��G��!��@-�H+�Y��5�!��`��[)ǫZ�qd4��GZ5l5�^��@6 A t1e���so�'�Y���L�p�_�������Ο<����}�	��v�nq��d.���J���lz~0�oӳ1�4<�uAծjx��Ԇ��������W�p������=.�Q�*�>6�:����L�]�ۚ����mt����*��?�1�tw�<$���Xk����JJ�*׿����ѫ�=AF`�X���5Fʭu@�E�yY�l`��䳪�b��cslY���P����d��^�C�\eED�{��6P�]������`���\�yA�|�-���y�r��yF��Mu�?̽�I �4�*'�y��������c �Gކ(\5j�8�p��ӕ���h��1F�)�Jc�/�C׶����=ho�K0�뷱�"�y؏�nߩ5�%~�b��Z-��%�6\��y������L��긖��x1�?�鉿�8�G<(`j��&nV�;����b���b��s�j�\�`���ٙ���y����F��HG1�g*K��������o��?�Axb̜�#��M�'�)��4-őR��2WGdP�x��#.�t�G "��au���VX�t����<�)}ѽ_�kAv�����h�FO�;�;�f��G�w�
����J�Ji�7	ח�o������b𰢔�R@��BJ��dh�]�o7��)�O���� �|S����;y=�43i
`!���1*���M�%>�&m�Af�'` ��+��D�>��H�ߟ}�Y�-IO��!�U+���c���zj`%�d�=�x�jPZs+�) $�4����n<aEMUS$c�y�o�������j_��UW#���2����8)P�H����ي��3�N��E[%M��z�nXa�S����;p�����Z��$c��V�O���>Rq��Kg�:~�������O��!w�"	.���K��u��+eүs���2^�@��6u�e�ĳ���kw���V���¥�'s&�{9�2��%Hט��Qx}�7�[0���
��MЯ� ����\�� R5��^��0����ؖ$�70����R8�H���aB���ˁ�����НK���"Ws����͌�_������[�Jze'�ݬM��}������$4!�Q��l5�t�~P��B>�d�8yl�e��V�+�$-������,]XJ����c�z�t�{wĵM�|�e��¤P���\���{Zc�o�%�(=T6=�B��8�G�E���mT��671C��Mℶ&܂�"���+0�>�5!e�H%������3峤�B-=�A�%`�s�r���/�H ��]������/�˖��f��a�j ���Z��+���b7%	����e1HS ,�(b��'Դ�	E�|�=4#6���rL��i��;o�������(`�4(�t#J�t7HHÐ

J7�����twI�"%9����}�����<�޳�^�z�s�	M۸ y���=$16=~�MD׹�Y��]\�������S���j����zO־&��������f,���knvT��S^xX@Oz���#
�8*?coɘ�(/�0;n��6�W�τ���v�`�Ӈ %��.!��(Z�5	U|���;�Ʃ�٘Fމ����8��O�od�[�)�}�s7�o��Xº��g���[V���wp�0��$�����ǺQX�ndf����'�뎖D�8���K������?�l|y��dV�-��9����g%��>:6��W]��E��M�ǋ��b�O�>}���t�����Z�-�@�U7Ǔ�s������?�/�/�H ^����Wy�qj�|a9�Ymi.�:F�����7�9�Q�^[ο�����*���~�,�S�O�cϷ^E�~�j8�S&�ix,I��E�DR6F����{R=*t_'�q�Y����@�n�V��I!���5|��ծ�X��RT��o��t���K=K�"n5Y�V�72vC�?��Me��D�\�lsS�͠����굄67�|����|��}�b�n�����aVo?}%��c&�Ocu�?��U�ң�p�;qͮZq1��Y[�HJ���w�����p�JZ9
���@��:uy��K�Ew�Lc�͎ֈ�
{kRa?�W����)��}]&Yx.T�����MjU��VE}}7u�n^��9�!�]�dhw@r�(u�q����3������l)�y*Ns��Z��&�7oD�k.��W=-UϤ����괚�uܔ@�`�-fxײ����&�S�*P���)$���z�]t� :�IF��W���s��Ȗ�6��V3��G/�h�t�y���J�_�
�8�@��d����������Ld��՗̸�n��+�CN5>��K�D>�1�������F�V�Ov��{�9�ƒ����$J�^�h$Ǹc�i+W��{�iB���u��Y��g*8�St�,Us�y)���m��4�c	���ӄ?�<J���_`Pz���ޟ��y���t(�-�=�˦5��p�ha
�U��3�����B���z�j�A�
ߎ��g^9�qCOf!LM}������Y����t�M��#C'�|�߸T^:�F,�3H:
����C,q<xL����y<DRۑ����$>{mHyܓ;��>D�y}r�=c�B��߿k�bF�:b0:����v��;��!Dd�_�3�<��|ˤ�T7�ζ�#~OI����><3y�\��O��~��-�tu��oؘ���7�̱̇v46�87{����~.d����]:�:6��◑����M�Ԇυ[�v�����*����2� �	�-����](Ƃ�ݹ�sڵ>���ޅy<���j9ӟ���&3v���H�)W�c��;j���k��[�x���`��7?c�`��>�����x�~�祪<��?��[��%�/�bz(������wދ#*����7���>���"y�ƫ�hTqM	�dx������j��$�dz��Ø�U�7/�=~��A\T�§������؟4	��I���&!��<6:
ݖ���1o��ߒ��Z��R���,�k��'D��`�t5>���;�c��:4�S0�>���?�'<�����F%&���c�+��Z�11��\�SX8�ӌ��}����͵�ۿ��|��M��}n��1M��H����[Ax�S���Z�.ZVN�YA�G�/y�1}uKu�'�n�=�LQ߆�E|qƉ��	N��PJ��e� y��=G��H]X:������6!�<�_���XaD]�8�i0��tr�l�թ�E��6���0�uU;��V�xU��'H���*�yu�rM�^�<��/�+_�U��;�lN�_T�J"MjC[�O�|h��V��V�uj�rde��[�UL�[Sk���	Y�2(�����SM"RA/m�#C�յ���ߏ���{1ʨ�R.%D��򨱨��O��xt|o=�+�Jɬ�wg���%ɖ�S���6�ʼ��[�+]�r[8�&��O���V1���Vʱ�D������Nq���*W��f{�z���z�y�A����A}2ns�3kYPGN�0�궜�Mmf;��*X��2+�#M�*f��Zg�X�o�0D
ON�c��5�f��ڇ?r��E	�b��k�>�cƽ�Űᓢ\�� -��Z�˂i��N������?����C*�u{r^��p�mw��;z�x�7X�>3�:���f�4��@d~����B]!�q�̷�)��
���Yo
#Xb��p[z�(dW�r'tn��oจ�бo]��x�۹�����},bJy��[߀�nhW����w.��cQz���|��Hc\�H��9%;���K��Ym�<Y�o׫��,@:��c9ť8^���<eT3T�~��kf�zm��,1`~��qۤ����I9�σ��*\��;�7O��V-�/��/�?x��2ʜ��_�b�?�����@<�U)ӽ��<YM���.��t�rk���3�O��q���`>�\r.96r�i��蘿24^S&7T.���XIt����Z��b�V������>��v>M��,�^�M/!*�'̖}�m�0_bM���YNG)~���Dc⇊�5����&J2�)�o�bN�{5�����I��_��9�?j���v��N �ش?�����$<e8@w���X������"�b�De��2H�9���b]��l��wF�[�A�"A�3.����F�C������W�/���&���M��c�����Q���tc2+ޘ��VHv�]�O8��]t�^���DR1w*��w�7��:+��Z���V��կ�;^[X��Z$X��Zl.����a��
���~gw��t&��M�~II9V�X���@O��#�
���}G������ˣ$�9������������To�>f��̧F#[c�~�"Ĝ�$.:E���F��x+�kSdh�?�FS��u���,�S�YՑ�G�Q��n�5���R��ݭ��fUcX^��|��w������cJ�࠶�=���t����.5N����JPQ4^�e�sȹZ��G3�)#U.ڑj�2"��l�,���ʱ�y-J�	6n�T��.��m��B�r����������v¬<���%�S�O�̱>�Wc���AE�wu��
Ε���Vy���o�ꝕRC�tcm��~����4����7#��88Ոn��JĠV}�p��
U0;�`}~�ũ��Q/f�d��01kc��G΂l��I&�b�{2��n[s����RS�����ɢ����<����B�_DwĐ��R;( )(�u�>�=i�N�4��O�x�2zu�d"+��b?�J�I��AlJR�A�t�2�>n}�LC��=�cU��h���$�De#���X\�p�P��M=���K��YZ��5��H���1:5��xd��2V_�m3mܶ�����:#�����.z�ZЏ�p�w��C��j��Xa�)�ʙN�fN�x��`�\]@�"�&�?챯���%1U��|D�EC[ڷ5"���<���ny��ȃ�==�H��ȣ��Ѩ%k4|�<��<�=��p�]��}��d.81���f͝���$���ܽ�i�U�a���t�[���F�9A�`���i���'�bv����m�!�7��p���{�덥��͹��,��8��8��sZڠ�?a�{�/�̌�Q�cQ�_�U�]��3��=s��ގ���6��%;�2��u�E�\�!��>�� ���Hht���F�Ռ��$�LD�:��?p��DF���ޛ�ټ��u��Qo��A5	�����݄GF2�����m��~���>�h�9mu����}q�i<u>���np·N�~��݋<O�H���v�v���Ѥu���.*So���q���پ&\��bT�r�&¶�(��u��[^>�D�t��	*-��]���9fl]�������������? m�T�v��M�sE�5�W��ۃ/U���3��ڧ<{y��Sf�3nPgUk;U���S���/�'<���?#N�p���w�m�ot�i���d��ݿ��|��㓆��{.nl�(���]�w)�Ջ�
�O�Rɔk F�%F)��8��s{�R�pI&�V�����y�7?�s�S� ���&�X����$�Hħ��ãN�;�y0��Ρ-��?�M���o&+~3S.�3�0��EX�70)>���Ly!$�천�O��i�Jt���<+��%��Ʃ0���$s��9	���`'C��q!�~�O;oE<����vև��B���U�\@�q&�jk�_X����5Xl�����|���,B 5�Nc�9nj�S� ��Ñ�r���fM��	���S��W\�P	�X��V"�v��7A+&:vc۽�{��g���uR���E�Kj< ��	֎�W�?��)�.t����o߂!�fE>Nm���'�K�����b��Ԯ}�^�R9�d�������Y�2��L=d���	C�I��l�AWO	��<���0�1�S{�������-�ӝr;I�$�!���p$i���y%4�,,����f���h��������a�Ɠy����Ӭ�d��`�Eo~���<ߟ�v�k?����Ie�\�;�i�l̞>e/e�̬!;���'U�T�SZE�OQ��E�'$�j���B�˟&Mn��0%G��w3W
�p��_M䈿�� �2�{�i�x��XI�WݤL�7�jؼ�xґ�%�	�V4�/��e�+%.���X|�(�#10vprZx�7?�'��6!!}W�l昉gG8M7�sҧ}��Y���%�R^�L���ۘmMs��e����ԾW��I5V��+������e�&�=�����Ц˟r������D^T���TGl�y���zk=���G?��p.��/�Bۼ�j�'�D�|�9�(M�w�����}��5�1͝ʪ��n\F'���=��=Sw����v��v�د]6�oy_�e�\��i����dWgd�L�C��u�wzZ!�'871�.����ӏc��%�jx�	��0���E6���*7�ׄ�*���'�*���YC�/�x8��~����/����53��(�Z��|P�M;U�uڦ��F'5��}��e�T���=��{�m��U�
��:/��	k����t��Wf����*�*�n��jze��I��佃��ťÏ���.�
h/�tf�LŹ�mf]�����B.-�@%6�7M�󤀜�Հk��ҩ��W���@���
0��ݴA"�z�6C���>��xW��0?}�$�}��ϛ�m�-N�	�(#x����a}6G(|�骓����ˤ&h�k8.�Ą�ݖ��l����ёYe�Uf�H;�����q����`�[ǊvJ�-:q�u0A�����^���cs3���~em	'e���i1l�G~8�9I�3�|�8�����s�f&���va#�/b�7�k�� !���{[=�(%1;;�磬� ��pT�1q�>���������@q.*Ӵ�ʣ�XS�l<�K�
����k���?�?v,e\Č/�J��������$��c�6g���&ҋu��7HxX���=鼾�|\b�<�KK�!��ǫ�(�1^����b��1LQ�Wg�xNwwu'e��ɼ���xp�|�=�����G��IV<���Cީ���+;�W�	��F�aL�U�����!�U��i�%��3��V����-�#��6~*��)�ͤ<�
-b�u�*a���mlb�nP�IE��z��H��,����4m�d����1����|+����a�G��������1�n�Z.��*y�%��Lԣ��K��Se(�P2�e�V�򠭦�]�)�����vx�w����lŐ�77mm5!O��G��k�R*��8mV�o��:��Z�Ʒ��&�,3����͏V�b�5�������Q�������Y��:����bu�����j#������H�a�����'N�o��|�qRT\�������M�m�(6��{mq�Q���+&��P��ׅ�#�
�ܸB�>��^�QD�ʯI)���`����}��{2����@	��.+;�lb���8M�R��C|yKZ�@��;�'��D��!A*hNi�m5�1.�e����D�T�u3�% �4 +AmKo>\T��mt��������?8�Q�ܭ����m��L�9���q|��`��������Q��r*�n1�{3^�L��Q�z�{}=�a����OV�[�!�^���@!r�Gf���$s��j^N�ջ,���e���OiB�x!�7��aU#�����r{�N�f��4εk
�R��*_��.�F�������q�VF��>�ݠ�7'+����;�ʙp,C+�S�!������p����|b*J����Q@���py�y3��U�r����o�a~�Y��C��G�pUk�JFH�V�{�4Ω���`
}������Ӟ��m�.3����������������E��tGT��b���c�	�F��o��b~m��3?���!N@�fl�z'���ډ(G�j�=C�9"�|B��q��?,�[/�zޤ!xA-��l�]��sX��K��i�hH�$uy
>%j�����'�^5�{o�,�Cb\C*�-��^�Q�aV��l�a���b��:����ޤ��q��:�2$G�Έf�|��?�U������d��&ۤ�S�;��w )��?���>G��s���7q,[���fēS't�����_=Q�#P��T�H��/XR�U�P"P��)��pn� ��7�.��\���5�ȹy�����Tp����5�E��qԛi5=c�m�b��T;|y�����suv5��v���'9�߫�)�)~�6��Lw���]R��omJh8��><I�,:j�4�=�dh�A�\�ݡ���g�~�]e��2�S���ÑA}�>,�vMv�H��
��(�sd�>��{��;��q~��l�f�W"��;�j�Dc���"3�/<6Y�w�)��ww{i�T<���_�L�\�~؀�o�^�B�1UcMv�N*�B�ٷ�t�2�+�a�
���"�u%1��U�89�{�����:-_�R�W��֭f�<��lU�8��"�6Ȼ��a~"�a�1�\�G��z "RY�Q����W��&���/���6�r���<�����$fH|�"4p��1���E�<���c{�q���˩��F�{7>U����w~}WSR;�S��vm�%#������<D2�N�c��S)+�0t�<�h��÷��t��ԠGx+���qa���44����B�X�:i�j�Χ��]��c�B��G7?�]��-�V���}�ʓ���I�	��1�����B?&۰�4�I�q�Po�6�:��٬���܃�I���/^D� ���dv�ګ�ȳ�uk�yI|Uq�35w؊�̌����[rF<�֡ǝ3V�s����>rrP���
N�#�2�uC������/>��O
��+��?5�7O�k:V*(�	]!wxp���~����"�6�lY�������`մ;^12��]�l<ˣ��(�Q�n�p��#������$Y�=,w���gj�^Z�9�kq�8c���0'5��cFg>���~|�\A�/Fه�CW��X��h}�̀�"8� ��:�O��ޘ��5�q;S����2�@g�9���oZ�����?���ˠƈ/eT�#�F��Ј�2/�[�4z'O�gZN�>��z�|v��w��y����D��҉xn-��5rf�f��#O��gc$"�q4�Y�i..{��zm��E�x�:ǥ$�+���]��!7����yq&(�Ԗ���S�Q'7�������*K����iFO�u�P���B}��}�w�Y��:E�?��7�z'�)1��&��{���p����Q-twůuz.�)ΰ�1�1�T	���k!���-M�	�6��tULh��H�7xT�%�1�j���x�Do~�YP��H�T��~|�r�n̬C�^�;�*gt���rZ�0�b3�������&�k�s'eU�{�54�{F\�Yq&}�����Ȼz5�*Ը�����mgt�ͧ�~��+���fB{S٘�h����{�T�`(!�#��a ��r�\_�b��Xsd�|�ag��ۑ2�VY0[���Y�z<UD��-5��[��U�j� �Ky��:�]
f�l���+�Mq�8��)�zK:r����?�O����wR9Bש^��}���l��)�Ã���P����|R�G��Km)E�4ך����ƥק���i�}��vW�-�=���"�>%��M��gC��������,���� $��pZ�KPA�9$M-'tV:T�#�>��ѝh!�(A?���Rx�}}|��'�B����)�:i�m��������2<���0��С�p�*煔��s�o�4��}Ǚ�+��q1��C:�g�)�o�]b:�*�\Jz���˿0��m�6Kbv'��b�F��;Ű����g����}Ey4ua�0�pY���ZԶ�ɛ;���Ib{�����ua)F�Y� �_9G��/����2H��C��ld���겉ͽ���2���5rN�L�QL�
��SL��j��y��5�y�V�s�+�����5-��8����?s��u�'�?�����X�J�S�NH;q��ؗ�t�{�Y���}�R_u?]�8᯷��$��K�]2�jB�`�U��+ .�wk,kvj�J�����i?@|EI5e�+?��Z4�ߟR�{�߸aFڿN���ڔ�����1?3$r�I���ה��]_����8Mv�,YN+��r���{��ɂã�EčYC�ۣ�.g��:�#��y��^���=��ܗ�Ñ���͈?�棯Te�dW��;�L�;�"�1�yL�'�_a��b��j�dN;��x�?,WN�]\�r�P���!ts��
��t�˭)�X�Y�'q���ً��e�+��n+g�z��(:�x�BT#x^�oc;��;wH��g�� }���Y���f<��~	�Ǆq�}��@��*��K���:;b�r�0�qq���Ͼ�S����>�sw�c��ɘS(<<��(E�����뽉�(����:���������~�k��K�OO��9�z�rJF�X	��������Ն��p��^����H袎��)��u/SK)�.�M�����*0+�t��"��,Mn��ɺC����WrΘ4�2����Y���:�U7I�2L�A�Q�a3��^���I_�mxʉ�KV	�� <r���ֶ�7f���4��B�3F�3�4�ē� �g�i�O38�D|#��	�V�6�>�����,<�$������ڿEJ�2��	2.��wgrhI���IQ�����Y_��cRE�L-)�mG�1�����6��m�/�����9��r7��z;�~�$���852^�Q�ԗ�����O^����-����ˌ���[h�� U��ZU�r��b�1��y��^��)��7$��~R���w{�GY}2_��~B�/8�4n,L�܎ߵ��4��u��a��8b(Qg?r�W�r�9����z�J%\��૮v���h��M�#���pz��E�9�6�J��N͠�8���,��:�ԕ�X
c"�0��B\V�4㆏�*y��^�5��N�_<�����:��څ�_(��ñ�"�K���'�z��g��Ky�BiEt{�����I��p��ҋק͔�	�'KbQ��/�]-F6t���jO�X���[��+�ũf>�&�G��ŔToB4OĴ+�f��ʒ�H���qDǙ�/��5�܌dw�:�M�:��*^-���1d�Nh���})�����y��t����Y�Gs�
a,d6#��_��-_X��Y<�{���sw>e[g��`S����%������������<r�P�2����C�}y:� �Y��*�]}�h�:�_�hT�i#p1�]�zw4��&m�7�������s
Tz�4�i��jǜa�`��bͪV�^V�Έ5Y}���:�b}?�a���.�yu��N�������%/�96)��)]ZШ\�&<�IЫU:���7���A�5=yS̧k����υ.��0+�j����f�ph�S.vcڇ
�t�D�+���N�o�l�ĺ�L>>��x��Y|��M�,��a�)�g���.�W-#��A܊��"���o\z�e��YO��;t�6�,�GFgyđ2���t�P�M����=��,j:1��{�LO���HZ��pqKȓ����4�=�����WF�ȆhJ9}�����9Ś���6�@�>�$���/�������0m���c�X����z�bA�|����#t��|�ĩ��kČWZWX��uA�'���ߓ��t�rs���g�>��]Я�cE�$�l8� LFW��_�NY��S����e�}�^e�=;�~����_ݼ�̫��8����t������F�:g<��.`��O�p����]��$N~�����ߡ�-��b��+��t������ڒ���e�UK{�Y���]s�g�����8���Й3<_��:l�xVYF�%��m�-tc�qŚ��9�I��.g^�ý�G�3e��"��P�*�&'�>��t�5�vίn��5���*nP-���ϼ���l6�^�� �E��E�v4�_N8�A�B�%�y"?�lը7kn�H͏�I'�6Fy�d��[?����c����K��(����=�U���c������5˧x#��I$���(Q�K�<���wl����ņ1�V�/cB����������n{	�B}�"�x��:���y����<�z�9�9�g֧�c����sT�I� �w')c�a-oe%�g��OF_�Zi|����gG��A|6���Æ�g����*s=x�2}[�	�{���E�|Uu�	����W�1�)c�9@=wb;�:ɭ ��Z/K���ǳ���D�#��r�N�����$�&��5�[������T���t�E��
#��9���b��#>�����q�>|B�)9�s��Y�5�!F���/V�U��~P8]�ిҩ
�]R �
a���z��W�L]���q���Rr0=����/�D�x�D~b�FS��	yK��m$�0��oؑp���ql's�(
�Z�6���k5�2�ۓ���/b��	<WR�P�oj,7���e�C�`��Ҙ*���,�� &'{����B����LYp�c��5rkh���_��0N4H��R%,��<z�EN�.�޶3ۯ�.�%e0��b&9.�8�d)���W�+�E��"���Xd��M��Ԉ� Y�g�Օ�\Q�C��MRv}��ի���>|J�[��es(I�ߵ�&_��+v��z�|�8��$$���m?ZkzR0����q�����T�-�uop�?�y6�4Qh%�� �yw��yI�>���a����t��ƀp�UH=7�P�a#?w�[Ӕ��y�̃GX|�sD�yʫ��)g";�Q�.�4�/5�w���)}�٬˥�Z�Q\Z8�ܨ�b�� (oH����oq�o׉J������e��?��8-T�>�S���P��n3k��H���͢�w�����j#6��?
��R�����<�9�'7uʽ����I��#S8��B�m���W�)Y��' <���������_^���l����B�G��|���F��o=�Mܪ���щ/LN��u���u����;��d�^���Xmm�z�;��^�t.�ը�m\:b4�r���z���޴�`��r��P��>w��ǡ�Ja�Ke$�pE��'�N�:}��"�]!{wQ���i��x3}	w+f���!��+C���T |B�7ڊq��I����K_�m�������y�ҁ���;�6jY.��C���i3���s�v&e��*�:��(�&�~�������R)N���rM�SX��:�~�'�qt�������Fc��5~��:�5_�������%����^<֯Ҹ;nW8�S+T�)�٬�?��y��q��g\Dw�#������;�b���]g���1s�̸GNgU��Ow�����>8��??sW�o�U��Y��d�J!�^��Y�O�?�b�4�g���6hls-��=}��Ӯ�?�̡򬞶�i������a'?=��|��@�~2Y���ϼA����O��tI�!�^+��soefn<�Y�����@��oV�bVIG3��w�V8�Y{Ud%
O�{�R7ҀX틴���m��$:�:#wx���4�i�Ġ%b�H[@�]���u�D�:�qjkp�hܸ9*�aщr�d�vtq( �w�R���X ���ɛ$�������.(m���B�:QQߴ��c}
:��o����k��s�1	��:ۃ��Gp�|���s�	ڭ_r�/
+����r
�V+��,�Q�mj�$�H�������W3�A���=�柃SI��'�uRw�mgS4j"E�8�9e!9,R#�'���������2ES/�T�%O����d�kz4BY��ri�aP��rpl&['qX�CW�K�����n[�|٭���=ʷ�˟��[��J�Y�l�'{�����6����ߡ
!V}Cr++����mBWt����J��#�2]6r;O;!G�(:EǛ��sOMM����b���5��g ���ܓ���fe��켘��'q�'��'�x�����5�;e�a3���ߋ����7�uI���ao[��Y�n�F�t=M���@^}���O_:QQlp@�s t;X��NЖt�����a ���ã�napsV��I����fł��+�fT�,�f�Px˒�#��)))�w&���@Gx��I��w�Z	�`�Fڒ�m�,0X.E�c��u�S7� b���:��yi��]Ip�}  ��Ȅ������#����\t�jb2��)�{�o��b*F ����+z�A
$D��db:�6�5%~�b��H��E<�?+D�EhI�PK���j��_���f�ڄ�m0XY1�>��k�7�u~��th0;��+�>�E�Y�<���� 
m]� �]�(���h���8�x����f�ԁ���]t� |iSh�'8������6"h�kPZ{�ԳX3���E��r���4+`uq�+���#hl�b<��5�i��GP7�n�o��]@��~�z�v�G��<�P�"'6y�9&����F� H?_���h�F ���`�⠇Qu)K ��Cv�
����J���*�����E�r��D����q��wP �_
��>t/�~�6�������z>��Xb��8x��Qy@ކ'B�3�{{E�D�A�gH��+h��dm�b���{9��=t�������2�r^l���5^:D߾
A!�=	����wB
��ǋ:L�3jї��z��C3((ͮ&f�6�� �H)����@��?��E�`�3�n4�@sL@���p�wL��4
�OB�Я��f���t���=�H�R0U�T��~!�G���)4��BHp5�r뷐��=� OBH~�P'������Ӳ�:Y���%(���@Pw|��4� �y�q��2	�,@J��0p�&��:�on��n��&�P��nyI2�%4D�D��`��A��Ac'h�K��F�Sh�$Wv�Cy��x��� �eL�� �����560P�!���"IVP�DZ�� ִ	^h6�-���!�w@�a�ڄ�Ҟ�(v��Ӣ*'|N݋Y�}"~���`� x�����x�Ā�*�֖~"������'Y�	 i2�^a���ꠜ4���6�������܇2��b
�R����: -�@9���,_8_h7H�?��,X
\c��H A�i����/A�^���m�א�p3�O�`�S	��fK0�EEm�#�����|��	���Y�O}k$�
v� *�*�7z�� �O��s^�r�훐D@��(���"�w�+�?�e���!Y%�6��i?�y��t����C�x�@�
��W�Et���@���!�	y���~��M�ߓ@��O���$=U��%շ$  �x�� P\7 a>��A��0��m�.�v �)��4{=��!��>W,{��6t2=��)�����Ø�����i�v@�P��ڵ'0�A{åe�A��~�*f�� �y��4���K��^Q�2�xC�M�@�������& �k�
��.� !��������?	]�xE!�ݡ]:�D
,��ܐ�w@rCDJJ��r�Ȳ	!�����@A�M�[' B��f+u�d0c3mB0?�^�8&/�H � �!�/�ԥ&B؃�:��8 �� ��%�X	�n� ��� P��ă�eL��ǐ�!�9@�(_�%�A��.)"BA��Ϟ`����	�/��&��, ��P�@����߃X|�����A���%ȋ��7c_y
p��+D� cȪ�mD����
����Â=ć�����4���C�S��j����0��20o=�|I�:q�P���2�?�&�!�K���C^@O�7��#�q��Z_͘L@������Rt�)���w�S!]gC���Ѿ�?��q��x�y-<����A����}������?���9{g��.ĕ	�z��N�$��! �2���{���O(���/QA��k~����7��,��ѐ ��x��J!k-~2�tl�ԃ�)D�� Fӂj�Ex���|' ���D�פ���m���4���q�W��xW�*��W�3У�����������m�s��B<�����FA�u�Ĕ ���֞
��W"�5�{xv������;Z^��$!�����**Am9A��֒�P���R�?kWu��讦�Ax�0�	��6ӿ�v��?B�����o�-����?k�� Y	A�F"��������]���j��7�i WX��'�/L�7�p ��m)�r���C7)��:���hf�\'W���2�7o(P&ea����i8�n�� �P�U��(5��ǂ�C��v�H$���AEf��MЍ�[Z�G��U|�� ��[����qKY0Y�'{`B㗼�Y�gP��_@��������	B��
�%�q��,3�L� =8/_y�U��R� �<C݀��~"*4Q�ԃ�0*77�|.6��@�����io�L[ �	Hwm}v�.E�&�h;�A�%M�r�	hI���������#ٟC|٠���bA�_��}�"�
�#��
���#"#-��a��W{'A���@�s;m<0ڪ�e*�d~*G2�*��|��Dx��ҭ�/���C��L����N�F�9\pa����m>�����vl�O���-�t����ꂜ�5К�Z�|u�ُg�6!k#6����0ns�@"����tV�jw �\U@؏_e�zq��|�j�����5)U�KѹN�a�EK{�^�oHF��`���&/��o���o@�ܘ��X��_=@x��N� 2Q [7�J����9|�!�	���1Q�aO�^tM�:��w�l�i�[��c{�*yi���Y ��L����Ś���	�l�����s��8�8_ FC�.C��A��7�	x�խԗ�|:�LC4ׯ�:FA�r���W�L�y@�����3T�S�j�fL�?��w�R�m�<�@�s�S�Q�CR���b�|i2�_=��}�����c��}p|	����7I����Y�h}M���\rY�UL�n?_��`s%���5�uG�Er�5��Y�Ů;e�$^�	����,S����})��-�v�,s�I=��r�ww�A=��S��<�㉚:4p����{��۔���C��8���. �P���K�%����_���n$��{�2D��՞����^C&�ٰF�ܸK0d�+�������־�kbj�1���,X�I�=|�3m�e��`�~ຟZ$��[Gи �pW[`��,��Cdu7�(:P�a�@�`�����J��&ހ4)0(�w�M�m©%kL@��X���q�D��.��.Wb�m���T.�i�M���Q� ^�HJ�5 ������������4l	8��$��&����Q�$����\\�X��� *�Y��^�=[�p�:�mL&��N��
�
{��q6`Nq�g��S��1u [F`���L� T�E���u0C�w��z�N{d�i�F�d�ζ1��״p֐����	�e�|�)�怙�}���z1@�-�a�:�O�JW��m�'�Sy��$�	 �a��J�`�@�lE����ӛxl�`���వ5t_���7S.�ӿ�����2�~�Zv$��_[;���H#O���5�
���F�Q��t�J��F1_���p�ƹw<���2�Y�Rptu�-��=r#��J�e�f$	R^��z8h�	�=(q�(�2W0�:t�|Z�������;�����[�p��h ��"�(��lU�2-�E)D� j�N/c�b��N�f����,�-ѹ�g�x����W����S]M�y�[�AS���)$����ZL~,�}+ځ+���Rϧ�sQ�&M6f��O�;��?xw`-�� ^�o�|������p��S �� ���O�ȧ6@�U5@�P����TS�"�:��u=�]�ÌRV���
sC��5� /�3Aڍ�CI5��剮��m,Y=��- %�Q���������~+�������J�>��U�S�W.��#2���dV-ߡ<�� �1H�Y:�����Z�s% �.��Y���	���S��ӫ�j�
F]#r��B���'�F#��.z�@�B�<�l��=��tg?:��X�����J ,]Ȧ?�g�wб��Ȣ��`�6Q��	���l�f��=C�}+�����s��b�(\�P�X�V2&KF���!�� ��P$< � e֖`e; �(5q���UT���8e*��2�$�hG�Do�@/�hd@�a�	�U% Pt�]�y�L��&1��b��i<��z,+u����ıxp`��N�f�i_��zK�R�F���!��ȼ\2C9L�M�(-�A���:33_�%�J�Ϡ�l3OF6>�2�9���W�EVϨ���_6Fv��%�|��M��O������g	� nzh#<F�r8w�y�T�@����`�8�q,�
p���n�g���d�	|)�,��o9}t����=��P���1A�ʎ�m��p�2A^�t� .[*���ã�-�o�fc�1�� �j4�)�y���K����ӐR�]b�Vv,8}�T��,��M�7���]�wd�$[ݝ�� �;���q�<��i�EW�jX�4�d��۠%��!q�@SfL�����7	^);\��tV�'��[� ��h��M�4GP:��H.�@�^Pm8J��m�SAh7�)���]�a0:iـ"G
�_`��{�P��k��;��J3�5
|	=�TM����{���B�_�D����1�E� ���1j�X{�� ��u���0=++�V��Z�G�!D$$�.�lF�j}����'�������-z6�"r""<��TE@MA��Х*Ujh!X	D�H� %ҥ��J��tz	!����y��w���~a>��k��������.�����=u:>�����P9�/{�/�������H�'(�fd����~�U�W9Nf& e̜�Eq?\��A�4Z��AY��NpyW�7@�Y�(�V�^ѻ�hۭ����W�d�W��*y��Ӌ�vBw�~��?�o4�]p\��~��k=m���;m��E�oB7 �5�;��a�P�iM�����Rƙ�}Y�}��p?>��?f�����}���GO�(a��ҏ�tL!w�3��k�C���s��%��.��~��W,�z�l]�6p]�"3�ޓ�MR��s�g��w�4^����.�O5��y24]�ew�򛣯b�����5"��˳�'�F���ye3OV��m|3;*Rv� GEcPo���f�o�YK�_d�
6T�=�L�n,��#5]ܱZ'���5s�e�]t#��o<�����(�X=�u��^)~Q,'m֖ܞ+�����Կ��"�����9��_
f�/���W��uco!�?}�ނk��5��q�g7ll��@a����~�X��W"~�e�:����])���'.w`�bl��e�CfKF�w��Ա�,��&iXI�n��V�ցƳ����-����8�g���k�Ѵ��֝e��?±ԽlZy[H�rł�Ty��ԏ����-�icWA疙����6�M�A5�-����8ʵ6�N	��T���Q^�!�*������	��5�:��%ո�o��m��#���>�Fپ?7��,��Zߵ���D2S�p�+Ip�`�S<���W��wl%u�y�{.��.բ����UTs�(�ӏ�6�>�����y�3�Я��4|�X澝W�jpƓ�!VVY�'��/Dv����^c��3�	���h���cđ�������#=���.<� �ϾPf�m�P�s��|����%s[�T�G�T�;*0w�*��}�E�ܤ�7J��O����M1ph=�%���2ܵ��Zͦ�����$<'�^6�
(�h\�uֳ{�Ύ���u�f��k][9�}$�P,4
6y�~���~���	?��=�i�C��彺�����gV?��B����`ۉ2�Klg�E�ۙ�I��!˵��.z���=�d�n/*��Zq26���yn:/'�)���/�h����s+�c�~�J�}�t����@ɦ�x)��^z`g��x��>���myp)'���-�\Ph�����n�iY���v�7I�z�z�Aή����9�v�B,W�u��Sf�e��)������֓;��M	��vl%C��ȶ(���9x�o&($���$G��Qs�H	�x!t:;>���']��no�Ԣ�g����q��H돿�`�g�[���5���	����#/�ΐt0�V��h��LSu�^U��ɧ��Y�&�o&��-n�������^���ow&�^y:�j:���g� �|�{�`��|%
[?τ�?���J��}t79��^��o��@��)��צ���R3ٰ�>o������v���5�5��V�M�g�E�(^�`?�fs�d��BM�>����J�����N&��?'�%4�Z�&߽���&��,�{�/�;u�(���"y���o���L�X(#9��M<���(�@�.�2\o�;��V��3�}��wo�qa�׎ɧC��;�
Se����"��n�!)��uX�nAخ��N��Ɲ�e�/���"���)�t$�nab�iߥ�u-���:�~��Wϕ�EY� n\p����6��CI�j��[EZ��W��m�:eL	���������[�T@P����#M
+g���pG"�C�n�����r��$-lK��Is��n��S�	����|h�*�� ֞��e-	�9u=[�қ��ָ�e��Ql���	��7E'@�A�}���Irg��O4%�m�Z#�0�0�~s�'�@������I�f�F'�_;L���������A�W]0Y��g2�Q��z�f�Wpt}��˾��~��8?��3ek�:�M1�mk��^���ēj�H�����DfS�a~����Ej��z�!��ֿh����3۾�O[�����\�$��I�w�ϰ\�]ȡM�:)���4�]��RO4a,B��tS�NB�l��.٬����u��JY��G5�99@6IG�������F`v'h�,�/��b30*��2�������q��  uC���k6/�'��.�nD��=>��{V0hǄ�O���o�M�=+J�b�s��!��.�x:�M/�ϾO %�..9h��9-m�s�,R��H�e�����Ue҂2V�4,\X	��ȆC<�	{)�&-��j�j�1� X��D�ӄEV�	&��|�q��?�[�˖���v�CJ	����.�7��e{�)y����W�k4/E���� ���1�Ra�n�1`[7�uH���B�����?
�X�y��'ekz��Db��8��Y�j%�h4�Lj�e�G�A�3�Í�Ċo|Q��%g��QŇ�]���v��|�9�~�.�+�	񞼭o���EVőV�����fOCNp��CA6�BOhը_A�K���]ޛb�����l�5Ͷͥj��8P�?�/V�(�`7��+f���bjU��3j��*:��x��3�!�Ch�_�]���tuS��Y�B�"F?>X��@���w����d[,U�6�Ű5rowT�{3�416������
$��?"�/��M]�SMU ��7��W�Z_��:�6�$ح͙�P�2�.�`5F�kc�"D�f�g3qK/Q'��K���8�i���OYL�޿���5�'���]3R�ʱ��"���u�<�~O�ˡf� �L}��&g6�E��'��ܯ��g�� b�'��!�~w�W�V�N�����
K?���������S��S��z��J�[&��-������\��p\���K���A#eф�6�� ���/[M>u{h󾻒��A
�q����d�&����7�zsvc�f������̇�|ďWB!��L�E���F���LZ9��������|��3�����ցF�!�X���Ev���(kz�?�p�C7-U���跈�?哊�i��.��G��$'�s|2ȩ-cb��+��I�؉@i������)#E�{tӜ��꡵`���sJ)W��j8)p��z��BKJ�A���.)?Q@^ƿG�lw�ԏ����$�D��A���P'������9��D7`�^���R��J{y[��]W9�-=jͱ�6��L3ģ��Xt�-�)1�买�rP���.ю��/���4�6���gT?KB��38��=�����f�����^�ʪ�#�u�' R�ە�,o�@���{���o*B;�}W.���~g�ν �Y0~�-f���o�nI��x��7=i��-���;A�(0���b0���6����!��7y�5��bY�3���;~T���F�q)���HI����ߪ鱃��� M�QRF��rl�硧�[���&T {��Gy�+g��*�M��4�$`4J#��t����)2G��@uT=����=Fb�(
���6�rȍ���О����*d�F�����T]>�`�ހ�߷��\d1@�H̺"��wv����q�$/95�����ҥzC��'އ�"����]U�,�6���mllx�����-5}�D"p�^��#�fC!z�����ۛTY5B�|�Uy�J�rx�ǻ�h�*���^�]oy� �8��Owz>f�1��H�+��Rv���f5"��PP��O�$k,�7���J4�#���t�0�"O�� no̶Ԡ�4S�7V��7�?��hOnz�t	/�Y.�ڼ�%��eG��:��R��[hG��̝g	�����/IS??��uj&�q����ݨ�al)5a]P<y�X*�3��P��ؐ[�,��EK��<�g�ע8�n,Ǖ}��׆�T} {������V��������s���|{j�C�+��Y8�yK�s�tdb�JSC�q�5��IT�Pa�+�2S�$���q�A��oU.�ox(��܍^����i��m֥��<���e�7��{�_n��5[�)������W~��
X�����H� �y��k������95���Ȭ[$�-~/ͻ�����),7;.��y�Ӻc�f+Ո�"�ګ��[����-n��4�!6a�Z��%���-�Zķg��I�UZ���
�#�'�`�4���m�{�F�ꁦΕ���v�f�������6놭䟁r��/�����n]����@;�pd*���Y��p�xcEP�ܗB§����r��IIė߼�C�Pn�PSmcP��Z�����H���E�9V�i���X�P�����5n���w�OZ�wQ��7\��h�?��T�e��{�����Y���l�&���D���xOT�s��#=��(�E��QeKֲ�7�e�z��k�� -l�Z�)����d�G���F����l�Gm~8��*o�i	�D���E������'�k�tA��m��+�mJ��V�-qtj�����*W�}�֦�wMz��V����#I�$�֟b��(߯��c���jڃ��Ô0��:������� �՝��𥧿�yj˄�id��p��4o,ՠD�$w*��e�ZÅ�[R�^6=����� ���1i�
у��Of�e挾d]��j�0	���}L?����u5s�����4�(p�\8���=sbw�J5CG���i�5�?�yE�@h����VGQ��[�x�(�Mw zZc-�H+�P�A2}�>n���͞���w�_�׽I�4D{ܬ�'�#�[��h>��E @�,�?E��h�6S~�KLW��~��-� ���+�>�X���&�+K�23*_8�^�|̚^ďy�O�40�Ԧ�WL�4]x\�S�+�o�O BG��֯�EWV�%�r�Vs_8p�s�
�2D�/Ab�cI�Vo������|��&'���l����oL���D6/.�8 A�L�	�dQ�g����������j��U�5��+�y��}����m��[��^}P�I��j�4V�k�O�˜?���H��r�J�t�4
��dL�7� � ��1�qX�I�Eb�4ba��`�RBp����*u�6�9��܅E�����M9���O���7�&�9L>ɮi��D�� m�_��j�;=�D�Y`�S�n�7�*�D9ʪq��UD6<Hx�/E$3��~�T� �I�� ��A:?�m�KM"k01rDϝ���N2C��櫵���V�P����	p&�~:c���o�w��^�z�.�ɠC��#��CC�&us���	e~}ZܢM�~���"����� �c$'��G�a��v.�&5���W:Ow3q�Ȧ��_��9��|ɖ���EmAҴU������9p�� a �6��t�gi�v��YkA�/� ���]��˂mD�����ѩ�K�1���B��ؐ���Cw��e����QČ�G&��L�v�o#L�����1l&�=>�e�²|���0��X�)-݉9��2O	g�g���`k�4:9�/���o?Z��.�ى�?W�̎c���m�W_�뾁8T����m3����p��ߪP�H=�L2Ra,-'�߾E�N������[T�x���6Ќ��	�m4� ��w6�
fx#n*Y�
F��?���Eao�;H�d�ƌW*��ƨ17��K_B~MكKb���%7���oM���?3��NP��U  Q�*`�mY�tbPpG�����Fvȑ�tҊ���J��8~�;I˖mِc��t	�Z[�C��ǨT��5ʞl���g ���Ƈ��o4��?_���΁:������K8�(ٟ��,�ְ C��M��Ma�a$)�Mq�c��C5�4�`�SD�0��$o�XR��LE�!-K�0���� ��8-}S���D`�<7�{�_|^�07Pd���C}70$AY�Ugn�Ӫv>K7��}+򷲁�"ן��4�Y��`ZY�vM��t�("��rm�ʪ{��rL���y��&� �5%o @R�ay� #�PS���mJ���P╣�Y��G�ݨ�?d��YǷ`p�:
��J��M% ��S�m����e�w�~��LX�^��̂���dtwoT�	�������Юj� �b��Y��"t�0]��9���W�1�O�ۊ����JlE���E̓j��n�:���CFf���s�l����N�`w���]��[o�e�)�<h���I��q�W)ᮢٰ��cUm��}��k�R� ��d9�]0�0�ψ�u#d��R��9�R3�ʬ�kVI����^�N��UHD;� ����hY�8p�U^�W�*��W����H����13�͍=3��t��F5���$(UıΨ|/�X&���x#tf+\{�ՠ�`�Y{F�l`o�!Ur�����M�Z���s��*�-I!ݠ��QH��7�U^M�6VzH2h��%��z4M�k'�qc{ ��MX{�W�y����*����J�Y�.&�׫g~��B-ا;*���8&-2���ƈ��u���d����u"���h֖�k1�D�5�G�^��Z|�7�#�x�NBm"�i�����Z~�|�-b�Gy?l�kV���d�)��հζ�Y�����O��$'�sE�eam�#|�κRLB�^�o+����8	����発|�R��[?�U�ڒfۙpTmVۙ�2ȱY��e�}jm�$���oj��s���$�(�\tIm��f�V=O��x{��@6.�1kvw�m7a= ��Aݏz~B5�9:��4�R���;L����H	�'3��Z�3��@`��nw�]%6��(����v�(�q���`,hg����aj���+W�����/��1R��;:W� �̶��
eJ�$�Ąt����m�X'��~�<,ʂ�}�yS@:L#^�[9q���kk>��g� ���)b͹#:�g�%m��Z���׻�B��|94Z��3>��5(��]��&ɣ����}��&�HӉ`/�߷7J���k��Zqi�	�� &�޵}��eU����nE4������:�a���pE�	� �d�6.��2z��A�v�R�Vy P?��"	����A�|��&�LM���2��0�U�O�\P,�X�| [;��-l{�������'`��s4�}7+�\ɋ@�\�ơ�)�h��x*(�Q�h�2X(���#�D�����t�'L��&��r})�b�Ru7\����so�F�<Xm�s�c՞�f�s��T2�Ǯ�@�dm{�<?(����0��:�H���	����@;t#@{�s3�C
W�:ՅH?0��$򈱕~z���p�h�0X|��u�a��;}���h	T�8�~�]a~���!!���,�xQ�yWS��Z�j��Q���,� ]�z�aro1B�yP��E�ao�?ӡ�����^�;����4�(�5^>0` �U�)�q�?|�r��oajX-��QR~T#X�NK!n�ƒ<�P�'K�є�0~7 �Տ�مEN�QH!�\��O[+�_~��.���
r]i�O]=q�D`��!�M>�s*�Z���l������&߳O�?پ|S/�	���ĺu�Z�e!j��(�u�f�7�Ȣ������D��)��o��F�o�+H��Q$;Ԟ�i.�Jt�nq�� �F��x�!��֔W� D������QU��?6گд#�5g�Awo(�.�X(��t 3�-s���ɥH�_=��)�ƞ��wk�շ��j~Am�2�~�9��}�s�'u��ʴ&���6��L�j�qД ��'�����P�4F���k���RN���D`�s��~�Քq[�UeJ:u喗��Qa��]�:���&?����t��N����ɒ� �<�:��!��p�Wғ�S�y�wv�0b~��^��tf�u��ztƐR��>�Y�Y�fy��4�_x�l3F�`@hӸ��wu0��>�����y�N�+�����o[�W�pvب�@�U������ȳ�e>=�%�
�Rw[7�N�4�>t�R#�e�,��E���,y<u�{��V���(�JR�<VdsM0?*���b'X`*C�����r�R�ό����Ӱ��1y�PaN���԰�'YY5U���}���1�iG�);b�wf�1#8Y�Eͥ ڙ~���C�x�n��{�J`냘 ��8��Gb�xErۉ����u����M�� sn	N4�:n���͹�Z�ʃY��EW�Vyz��f�_ 8�R&K^��\~� �LC
�x%��7�{����ɚdk;�Ք~	��Q�SE&֩A����>;��Cx�L�#�?��43 ��9?�& �_����gbŌ����>�Za0i43��䮂R?R[�]�r��[Ul-"Mc�V'!�S#"f�X��W���r_{��D��Oޓ�:W["�)����5趲/�-.f�a�U�y�5xrD��@A�#Y���?y"J�#����\P�Poɪ�7�>@Ǖ�M��Zbn<7�5������
3�����qH~�ƭ�k%fw��u�8�~�E�/�.�� Tď�),X�*�ݑ�۵�(��w�o�pW{FƱ��� e�ƞ���M��(�x�+7��I�
�Xۜ=a�S�w�w��$0arR<T�nC6O;�"5��C馛�*����F�}�Խ�bZԣ�Cյ�)Yl��k`/���dq�7��>0���> h�#����M��F҃..�p�����=�XU�����d������ lo~��6I Z�1�2Ӟ�=}|uv[o��j�y:���HM�U<).��Z�s&��	::�x�~`�>��|���00`oW�+j��P�����N���kePM�`���u�{�a�_U��4��mϏy ��Dhd�fط�s&��`wҲ���_�ح� .  @ ��Z���9�SY�麄H5�\\�u�gf���V�E��ؕ�ULn�3ۤ��1�V@�U�K��m�L~����@�p1:�Z��J�=�'-X&C�+L1�K�������a�z�~5
�����E�4�)��T�Ct����geVʋ�j�J�>HO-Ϟ��n��ܬ��x\�J�����H$U�̓�����>�r����[xjmQ�� 8@�*�h�
(m@g���jһ�+Y �e�OjGdrb��,c�]���M�[m@�]-�����#����(*=�,= (��XFJ(�Y�Q�9��}>7�	0�s.���؜���I�;�!˓���G�k��C��E�ڛ�O#�w���D*#xJ��1S�K�)OM�9͝�~[�z�cfߞ��k�qvP�����0��̨�T>��zd|� ���T�wv<,�b�=<�U�ph�u&���i(2�h�%�D�2K��7�����!�WXF�l9'a�r�͑vy��rL���bc���|b�	�q2C X�
���`�ʦu��T����i{�������$n&���sc��̀>��X�hS�8��(�L�[��W���H�g~�KB(������˻�Ӽ��6�E�~	l��&"�H�{�B�1�LݼzRWM��əFȲ[6�Z���fW����+@QE���"'��D1��c#\h{C0���?����'��@����EU�P�A�ĭ�'7����mx�dFGR#��6�+�}�-��1�ǘH=><��A�T׭(���cyӉ.0�ת�a�&>�,�����ۛxt�5f��Td�p��=(�rS��c�T�J&���[�HM��$��s���?WpLҫo��D��)�fˍ	!����l���^v��MTg��!c%�a�AJ�jO� 	��o�R�԰��ⵙO?�(~�/!3`Y}�� 'S.�*F�&yZ{_Y.��G�J���Y���=oY���2����'��{~Z�yS�{`V#��-�Y��"sn�&��G�S��6 ���<3N͆�v @��k��obůtЧ5��!�v���#;4� ���ß ϕk��q����d����s�;���M��A��<(�h�[85k|���1�}����*��k�)��jF��m/1����FYA�K%�����So&f f'�a���gҹ&�V[�4����Y�SI ���������C�l��xo��jb�^��V�+��y����2FN`JV��^O#�#��Y�!b� t�o`�����>k&|���1x�א;`y����b�$o��]fc��<�s���Yj$�4|ߕ��r�/.pTO]�M�/�a13}�M�a}�k�0ݏ+�{Z��[�Ӆ��CK��Ͳ&��"�N ����d&Mւj�Ԓ)<��͂��ՇK��_�QTZ�4���^i�aL,��|W���,������ H-��b� ���c��KwʏsJ��e����*��~�1���i=(V�}/fϏxE!\�����r�{�"�+/��N�%4H��x���Е�V������F*&x��m��b_Uw�OGv�ږC��VV2ˑ�>m;�(|#9\��A��kJ*��j�0UA�$�h�?�
�1풐f����#͸�g�)k���<�?��D�q�ӞC�#Uբ�1���*����=Wf�*g�[R i�9��S���%��� �[����WI�����z�3����Q���7;�K՛�u�<;�����̂G���ɚ���e�_K�K�Ʒɥ��|	=|fu[��%*q�P6��n��l |���U�Q��2ﲇL��I�lwF@�M(��5~vVm��]S��S����_g} Rg�j�;+C܃F�V��qo�w�e�F��L��B�|uN���g7#H	��  aT,,dw��p�|�PB�M�M�9��pIh7��I�F���/ ��w 8�ʊ�f�H|x2P��*%*2j:r!�4��d�4�$��Yj%��.�~)�&CI���7����k)%���5������~�w��^�����8�W�90�R�]��3s�9��=��fl²��w�cfR���F��s��k�j}R||c/���U6(�2O<H���}��n~�CYI=��h��Z8J_�Kj�'Ƨ^<�$�����0�Ң���)�8�K��[>{��<�ln,���yR��K��Cϒka<�P��d�u�<R�D��O���[��h]Y~�u?]8]��	������f����QR��⚨��a~ڇ��w��Z��brI��S�\"�n1B�����
��ky �~X0vƬ:����ڻr��L�x�+(ͻ���
���״����ghl�Ҷ����=�,=�+&�Q��,�r{�D1�iLoi�lʐ�(qݮZ��T�1�����ni&�{Y�#���2ն���| ���K���݆^Aȥ3�3��
�su"~zN�ZLE��{�E.��f���X��K�;��=�/2po���v=����s����CЋ�;��ܽ,�*����~恮�,�-/��s���k_U:O&O����/�|�sa���v��G��Y-��7��0?B���a�C�:vH>�(u��[�����ۥ����u���j��߰��bP&��s�<���oWI�T�<$�����h�8�Rּ�畻�b�����L�t�:��_�$�T��3̟/m޿�@����&��!�[Ԥ�I���_Ȕf������۔�Es�ci\���j���J�zS�����O˲ ��'8��Q1ٓr����� �^�]|^9�ss(���n}Z��*��r_RCd[�.ޣ�̳W"�J��_3;;%��:��fI���鰍��@9�D"F
o
�e���|8k]��].����)PtKI�A�C�9p���d.��ioN�I�����Ç2����6��o�VQF(�]��zU[}�}��m쉣Y������s���S���j���YD#oT�Jg��l���*���4��%5U1����)� �˾x"�b�DGߕ�.#���n2@J���â6�f��Deg;!�������x����WE��/p�{��)q*O�o�Z�}h�P��4����O��Lƛ����	N�u�Mk]���G�ĩ��m���X��@n�Xմuv}/�A��� A�}E�lg�:��h�Y�_g���2�9���lWP,�"����v
���=
����Kg�������j��]M��	H���a����mCu��4\f�<%v�f�9ծj��>�#E�Tw��?-褤��_�������������yc��J�7�;��Vx��J�f~JhH���_��6�s.vӁw���4�I���y7JMw�R��u  QVg�.������`�G�U�n�����e���c;���_�n0ߟ�Ϭл1'qR'e�dTW���nT������K��kx��oU��qB�x�KY�2�E������N�,S̵ت�C蔏'A1�NƛS�:��a�\;V �5��±�YFl*�����{����2�/�DmhP
���I�,�y�ª�*�`o>-��~�#l�t�Hd��RX_ݕ�K��U���3�2�ʌv-6D��||:R��͋68'}eK�P�+z>�uCB�G"��-��:��Œ�!R�boK@6k�� �ݾ3�~W>��e��Y����2�#��a���`p��'�$k�dɷ�v�-d��k������|��l߿���o�'�ϱ���Y<�S�K�^���׉s���S�W��ߔ���X�@����}>��DX�
�u�TS'�m��6����B���f��[�ٮ1_��=����7,�<�zi�}aM��b�=�k�[~���}�� �:�>y/�������*h�,��!9heh�{J����7Ko~���Q��/9,�F�#��>��i�dz��vc�٤�⥃k\��ϏL�ǖ��1ȘYK}fR��5�����G�}⭆��J�	J�0��*F�}�����n0���Ȥ��KM콢mKC�C�T��J��ڬ���|W̫�m����δ{|Ot89� ��Z\H����)Y|,���l��d@�͝M�(jŒ9��i�'��.{_og$�ta���c�׬���݈��Abe���g�W'�����S�Z���	��"���-s?u�"�e�f��s�ՈOj7�i��NTF��-UL����ї�.��s����;E5nl1w� �F���[��a�����RK/m3'���f��� �)�UtUw���=�C�9j?�Fy�\{�_��N=�$`�@��h������>OВ�E���+Ay��a���&�2o
	�p�	��I����R��?��������.����g9[��]�v�d�[��n��A�#E\����|�}~50gQ�xnq!�P�B��䘿��sP��p%�dGM���h��y�9�3��j+ȶKJ1�Ė*��J��Mp@��p)x�I��Ĩ��s�b��\Z"�fӛ!�cja�ףЊ���ǘ��jwY�Bu���
3�+>r�������8m��B�z^Lg�Y�wߙ��vE7a�E�'p/��<~=d�
+�Z
�
��}<8��ԉE��#\�h{aD>�$usz�ٷ�v7�����_�U�ӷח�^����K
��+���.`;}�*�pB�U�BPø����m�
�S[��3�P\��H�?�n��3�T��z���Z�^��o�p�n�/�ϓ��I��^Ξ䎾�|~�����&���XEX���Wu8��)���wR��W=������330ҫ�R�Ng67����m<�y-z~�`�H���dS��,J�t�su�V>x��h���jn�x�rA�����C﷥���zw�W,�"|ld��_�6��]�2��fg�2g���0\&�zU�*�SY>�&;���q��T�S��3�w]U ��iͻ��.��c;,�����ZT$lpKT�_����_��8[�Z�wd7.�<=����D���dޅ���B�?`|%�%�F��P̑�<6�յ�~BJ�b,���D
��";:=���K�#p��DjQ]��g�_��v�	�C�j�>#�g��u��澋�$W��x�vZ��Nԓ���c������t�� �`Q����ߺ
��^dW?��S1��;�=�@��_�g����i��%6'�p�ؿ�R����S�-�� �~^�q�r�f�d�Ns�9qG�У���Dx���Z�����PK   }�X�F��^ ~% /   images/b0a0d881-65db-4735-bc7e-86e9309b8843.png�c�&A�-<m��m۶{ښ�m۶msڶu����m�x�s���o�Q���b�{�ZU�"�%`q`��� �KL�������!��L.oG�{�8+K�����;��臔��o���vSU׫�Z����e�gT���Q�J�(��	���z�1��FW�l�hYWe
/��%����lF�$�U�QV�?~���[O�[�Q���O�3ƚ���=��3��̣x�tpo��)����B0��儁�B0T ��� �� �����BB��J�������R2	@&W����?��Z�� �c!+
K-�YQx��?8���dg��	����?8L��g��������?8X`�4'�L�<��	���?81  ?�3����o� ?]t���3 ��%[�(�°�� ���_����_����_����_�������{{�gp܉y�%i��y������s��Ԭ�\u����\c-���{u{��礡�*}�K�M���}���tEA�{����=������`��]����c�VC���^��^.�]z1���6�n[k�Ս�`�է�S"ѻ��m�nZ���(I����$�w�Nz�zNDn�����>{c�	�&�띕�l'�cE$�`��Kڕ�Y�L�)�ܭ��!��BD�G��ٙ�Y�k���6%�턕���\�q�J|��F�/���]:%߅�i�4�pb߮\��|��=��@Ҋ~H�:�O�� �_������>�\h�u���#����c��kK���!�㾮~��@[\�5>x�$T�0���۹���3.�������o��}��u�S5����G��o�Џ�8����H^�H�wc���q�9L;�i��q��@g�s�%T��{mjq�����V�f��YKs� S(�t{B�nA��B4�Jݺ�|�m!Wss;��� K���JK���&jY	Cv[����E#�((��N#�6ٺF٘R�h��a�QCh����Fng�y�<\�����ե�@�*�l�-����7�J�.�>;���4uX��q�bK±������ �(W��,ʳ2Ҹ�ЈJy^�������F�z���5��vT���N7���Ca�*���Т��&@&��J���xc�`4>��8�ĵ�|�M���}t}�+�A���_M ���(���t.������m��e��d��׈�<��}��ݘI^��ʸ�
�1U3����,��4���B�c��y�gZ�y5k�<�?���d��`����ުB�89�5ٚ;��j��j�IҪ㩶*��]�,�S���?y�H�,���9n�����o�a�]�,��vm�[�k�ɡ�4.�A�c,��Yj�=�`9�����Jk|\v3�2;�d3�1��s�V��;��f���`���5����4��A�J���{�ӿFHQ�:i��m}a����������7�^ɔv�=m���,s�ai�2��<��-��Ai���~����La���D��������� h̹��&:���
�G�x�5^rv5�[�Z�0���/g> }�kh��V֌ס?[��;
/�B]-�[׫���gwa�<��1Tmz*F5�0߃�a��tዣfZ�q�ԉ8�T�u�:xk^�/c,f\>T`�����j�_3��RaK�r*�����+
�3�������W��F%,�i�� K�I�$���#O�T&:�F�|]��s�s���z���}���F�u7�HN|8�<Rz�=>ɚ%X��m�rN1��WP`( �9BD���ҥ	��X�8�d`��j;T �=n
s�w�ҙ!�� �]�<�J�۠�^�0ɡ�K%=��! �!��q3��M$�F�7<��"�"g8��{X@��)�5�ꤘ%2X9+1=�H�"w)�$��;�X+��Xc�)j=���S9H�^���bɛ�7YsX��s�$,s4�Ya�����l��l�r�d��!�tb����T̝��I~
��"��gV;]o%jU° ]e��,�'��I�'P��L�2ѧ�d����ݍcx�)��ڦ�k���6�Ü�����Fw�}Kg�@w��F��c�af��Fk2��j�W��0"�+��M���y��ƭA����_ޱ�ҿ���<�*=��&@�Kh�6�i*g����n��F@}����e��D�lb�g�u1�j���Nl�Y�bL���'�I��O��q��0��8��Ũ��N{�c��kw���2���b���j�����پ@ޡ֪:1R5��]����.F�L�7�?�E@����:��5�"��w��"�Atj�}���}��l%?���/m���L#wK���i}��k�������U��`(i�~�"��;:>�i.�<�QO��� ���������M��{�)��������=��)��w�T����#�Z��Tt��Lq��JZ�����:_uVB�;k�͇V�@	=���5��߃A|��*h�z5�PH\��A]�Q��\��c�v���X��Z詞i�C��i�v�G��5��<[�J#=ZhjvcFF���V��̣�����گ�~!��]MKo���ua��6�'��󸑈q#l�jM�y�`����8Q[�{�r���#]����j��0�ps5�̯&py�y���=��-��$y�نL��+Q<��Ů�@�W���qM)��^OX�����K�Q�����2�ʇ1�X�j]3s�:5,,�����r�'-fmA��S,��Ns�/ؘ�_�N��M����N
s�d�Eᑉ�������@�hڍ�h�)w�����leڵ�I�6d/Ժ\pI3�JULcL؟j�t-�̠��}tt�/�cia�ɣ�u�����?zq m0����b;s�3僗,i�|�I����8���,�d2Ƿ��\�Hqc
h�a)��]OA}ˮ�Ȣ��D��aD7�Iחu�jx�� ��Ϥ|1Ab��1l�������c'�]�;���N�+Z1�d�M0�cN�g�2�ʸ�Xͨ����J}�[�8z�5���:���vD�f���Xj��uml���ű�{<�����y�c-w��=�"<���U��M5��-�j���V[!D�9#<�=��n
Y������_W�βV�u7�Q6��������y��u�נq��ş��VTƐ!\F)CG�}��R*j�0��9�=�tU�j]�0N3����@����Dܱ�4q�-<�/*\��9���p�W|���	��L���^Ҧ�/$g��RU�������b�����n#u��6'h\�c��������/W�-���[S�T����=��J�[��g���IJmL��������J|筄>�*��C������=�$�}e�����A���l3D/���pm�2�@�˒\�(��d�o���W�����TY!���K!2����i8��V�?�'�f�.����&���������J�̙MF��Y�r��U�I
�S����đ$;xOr?/3����a�$! r%�X����]|����7Njw���(|,R��i�-@�u�༌��h��'�����%mF6+�&��S:8��ư*���a0^��~X�݌����κ�'&��G1�c-c@:��NT~,&M����?x�!-��\ә�u�e̲J�8&Rt��p`��8Q�b�n]�\qU-Id�[duv��V^5�jU�֎zdC%u��;��%��������$c�`U˗֧=�0���j����Ȍ�Oc�@ ��bf<@�Dg����.���W{%��0�`q���4%7	��RO�`i��Aj�l�$���%B� �-X�)���)���"��c�^c�u㊣�"
0�UF�	-ۆ���gm���֛[�niߥ�������H4�
U�& -�����p�Fef^&W�כHZ����N��$U�N�%[�y���]6R߆�r��N��rp�1>�o�����P�����O�2?V�����9Bu�˜,�;��Q��<&���/
�W�0սH���]�V2"�� �jkl� ���-{yY�I�!��񹪠�l5�X};ʈ#Ixqh�]��{����K���Ŀ�VM��ik�)�Wx$i!�l��`���yx�+I<M"ΔX�!:�=����ь+;/Pθd}v$�;Jٓ���^5CS�D��%U �����rj��k�ь�H������7@.^��N��x[��3������у�n�=��H���>���򣗿��ǿՆ3=�]�t�5�v�Ց~�HZ�(Qe��<+eY��~F��F$�b��y���^X���|��;7�XR���h߭["���P��0eA��f|:QɎo�U��o�
�����Bq�\u�>�j

�v_?���T��4X�p������������jVN��E5�>�%��g�Wm8L��N70�j`���}��.���;�(ԉe��5�^�)��	B��6�Nۍ�;�D)�<n����z�^��"�`� ��I^M��q�'�����T�ixq�'�\f�9n�0�ݔHE��Dμ,9�LBy�F	������,��a*��cMM�ʖ��О����Me�F�����8�PO�NQ{�A]>_,�����q�1б9��=��M$c������y��yX�K�XPl5g[����}C'�}�z�;��R��D��b4��B(��C���1!:�ٞ<RL�b�+ �����g�3��
��f?�W�燈
����:z�[}�(�O#K�T�I��^����5#t�	�i�U�y��he^���\t4�P�����f���qa�Aꊵ�%���>�ߦn_4�%|�e�-YLH�@e�h�,A�3z�=�`��eÿ7��P�+��EOڦ��V����i�Θƕ����p�{�eB�?��J���A�^\hq�����Ε�E���Ȣk��NYi��͇�b�舼HB��N"�Ob������t�}/V��+7�R������l ��"F\�B���JU��*���r�W㎑��T�D�P7�M;Li���H�	 ��F�nlL����Җ��t�$,������(f)� :�$!�YCceE��
��!m#1�:��2�q��"6���-�	Tʒ��N�.��7����J���a�yC�+ ��$�U�Bzϟ< 46�
ߏ� �Iw�����ǃI�b���_�m����=���o�Al�F$7����ܐP�N�*�yc:��w�������=�Ut��L����&f�B:?����U�B����?<����RMo�t0㨑���n�w���hB�1E�)�>��a�8�:B���Bm`8~>�?�^�)���(�0��������r��k����S���NW��K����~?/�o�M%V��~��N6l��y}�|I2�ٶ녤�)��݁z!8f��8��`��HG����+���C��0Ɵ�%P�{�A	zWI���q�xG�����$�Z�C(1�E��>T����+�L=�3�$:�ZF��yq�%�pQ�^Vm�"�D���t�����&(^�m�"���4\XⓉ�F�i���.V��(�����%�?T��ww�gc;%�`�w�/��3S.�����*R����a��a�_�r[��x���#OX�p����t��v�:4���u��W0�F��IU�^�rwج)N��4��C��m+�Z��U���C`�GZ�N^2�D3�)@﨧 �m(	ˬ.%�&�^7"�V�9���¦�����C?��f<���1|w���@Z��Sv�
(F�%DN�䒬��j�4�6M�ﱐ��տ�����M8��d�����W�
3�_�"M��1w/�� y8��J����aq�HQTq��ɓ�H��g�¡�͉�Oǚg<8��Y����L�#�B�P�(�����DUh�k;��4%ҳ%� 	ó��M�� u;���G/N�1������?� %;��J��c��;YK���=�J��p͛��!��V�~<�*[�O�����
_��=H����/��{2��$5�yd�Qz��
y��5Q&n�N�ΰ���Bc�����d��V~@�����>�|����2V�k������*#1�(��K�_���v��ԛBʱG��{����2&��z�������oz��qf�҄��P,�`��1��Gxt��Q*��?�J��*־�B��S L"��I|9y6N9�������[��78����@pD�.�-�
)ؙ^��i1A�%�ܧx|\*���3~�v�L���>�!B��G (=$E,h��~~��dD�9Q�2���D�� �;L���nYR�Md3�D�#+8�n,7F:(�Y��I��!�˝R3����ϓ�r������j�����r�?L��梵"�ˌ4b�聹���I Z�1��H�պ��eYiY{��{��h.p;�����ﷃ��T=8FQ''a&�n�e0�,Ck���b�[B��c�ם��췭�p=�.Zs�O�t0��,<�mJG�>~�|�5k"5[b�X�D��M/tR�Ħ\�Wb"��L��o�d^Jv'��MJ9���V��s?�����u�Q�6@�H�����lL>�ȶ�q����j0�S;̻a�t��M�7Y�[`p�|�Sv~W%x������J�����5��ZrIƋ-��0���S9&e�y<O���l��D>���`�JM�r�2��_���kVP��	^���M��ى�a{�nv�s#|��=ad�Q876�%P*u��������!g;Cw|��ؖ|�ļy���u���Tʈ�4�X��=)vϖ�Ռc 2Ѝ��L��y,)�qG<�A�����!�D~o�8����#��|�?,1
��ei\!&l4va�P�a���r�󁲨�D��'}Y�߿����r��S\�ӝ���r��H��:�Rz�4�t��?����w��f�J�z���ō��|�ZÓ�^�����i�6!?�BmI�d#@n.��n7�x��W��~�10)@q�ݣ��a2�H���n	�������-6�hM9�tC2%�dR��sh)2K�M1��;���QXZ��~uYۏ �������C��='�q�I�Њ,���J.= �] �Ϗ޽�8:BT%�X	R�ic����!�R��t,��R�y�a���]��T{��g#j����~��e?;�Ni���a�8��`E�E�����G�)��k��{s��ٕ�����~�J'���0��4;y*c�ջ�_~��S8�D���/b��x���R�
='k�k �9W@��L�865���(_�3'������$�0�����	��,<	̆����N�q$k2Z�0ngA�U��l|��MnεR�ı�f36�Y17�
S�����9�n���Tz6#0�-�}(�i�jjH��ˉ�K^-�<QQ-�R���D���VLH�JW�DN���
�O���?Z�U9<��l�v�W�+6%����`�ֆ��[�U����X�^XW1z��Ɖ�D������ ��dJ�y���ƱC٫u�0�������_�I:u�1}gxC�����]n�\"@ɶ��SN�UQ^7��fn^jG1s��}��*&b�	��כ!xt��l�Ê��3�� ����6sK�ң-p�z�ч�H;>律�eZ򸔶Y�֌\���e7�����y��b�����t=�u8~�������X��0fYT����Ѫ�W���������@���` ��,s�a�V�ftR?�q������̞?�{H`Ø2�n�9������Z7T�}IS�{H��F���n��,��~|U,����@�棊k�(jϵ#,@��*~�ք4�8 ��T�MZ�2��f!.�A� "0ه�NR�~��/&_� �i\x�K���
yV8H�2���ޯ����b��߽+����aXĳ���cT0p�����nSIJ7nDx��W��M�]s��v�ؒ�.���G�N�����,U!��Yss�ǭӖ�D��-�4�v]*'�UMĞ�^�o���4h��+��^�Nn��^g�� i�˭�sc)=�}�
��	��Q��L��m�@?��Y8=������E������%������y���y;��<cM��n���(�QL�1F��K&~��6ؙ��!D'����tE�9&�4dOיYz}������_;��ӛ�J;���naj����8� �V�a�����u��?dA�'Ù�\�uX�>]�9��Ű��gc�}ZI]�(�(d��F��{��']i}�MB#q�����-�,��Y�2�]F*e�B��(���j��L�9�Dv�U3��[�B���l���*;b�b���k����ʂm�� ���0!�.Z��f���?���z������%�Y,��\�A�1yt���fo�F�#+E���c�I���y,�0�F�Q\��o�|�E2�sH?�|٠���p� ��SO�9�{"�х,�;{�·��E��ęK��%����kT�JU�ݏ�u�Mg}o�}#C�v�_��_�3��&��_�������Q��n�x!�+ӟ�p��u|	?���n�q�z_M�z���q�Ǎ����7�"���}]gz���5��TRQ.Ө=��י6�s ��2����8��Ke���g��2 ՜Oz�9#����;�ҫ���ޗ��%
Y�-\��A4����T[��)OMR?���>z���f��c�;� �t���H6#,T�/T�7�o8�]�y����t����8b>x4�dQ�ɰ�h�+�Zrj}�/�D�`L7�H���+aj��A�j�5w5��P1���E���-9x_#e��k6�3�!����n�tD�{܁����~�ݍ&���3��q�\?��^�wm������(�z�Q���
��ד�M�ש!��� �/A�ƾ�ɤ&~����C�	�(3�̪I��%s���4.�� ��$\3&�)Z��F�8HY�l�^4��13���5���R}]���"���/�Њ���Z<�yw�K�hHPy��2�HN�\�ш��[�:�>ȵҏȼ��Ԫ:�L�u$�����E�S�]h ��51D�{��#W)�Vqא��{S�L[_z����!�*éV�B9{z����4|C������,�'�����&���Iy�'CZ�۵n��&�Z��*���sQ�0Kʽ�&�Ï^\�hVp;����Q�ԅ!<�[�++H�ߒ��{�Z����%�ȟ�m���gI\c��Ӹw�����*h*�_'�'��N���d����T�@fm	�c�l�
i��D��$PoG�)2�\С
X�D�PZ��j��l�*
2�F<�ͩQy��Y'�E9LW��P�eN��WL�0{\�i����C����lB���̻<��	�۵l�����X��0]�0����0����CG�R�Cw%v��c)P�=�ݻ�p7H}�3���_`/��/�<R?ag�	�hG"78��?���o%퇋.��>5���o�	����S~1G�9!��;K	��;F8���B84�b K�q�by��ie4 �����'5�&6��õx��^��Ȥ�$H�);f,߯��%�q�׷G2�\Ɏ���f	SB����m:m�j``��S���]E'8�N���l���>fK�LR��iŎM�a˓(�e�ŀ�y���΁���c���s~N�g���E�Rʋ��/n\�LDEc�_��v���$�Q ��P��YI���	�]���`�LF�Os�X_��[�u}�NE�ϕ����ߺ.΀�0@��A������ΟW�tD��tA74y�W��+��f�-\ѽS��+oD��	��z˹�ʙ�<���~��7����-a�z�(�2�z�;��v�&F��߅�~m�K[ʳ����2�ɵd��R�系y�L~��ܩ~� aN[T�J�����vk����<Z��L�͸��ͳ@��&9��WR.�P^���E���@Q����̓bt���'�
�k0�u�o!ի������!���g�u�������ym],qV�����UU�������z?�Vi�8<`��N֢��D�I��,��k��B����t/���^�I���\G�h(�(y~o�d�Z����$�]�1�1�x�@�9K�Ҥ#]A�e�@1E�Q3�pd��t��'y��.��&]��gS��~:v�j"@��"'~��Ŗ^s���.�j�!}m���M��`<�_�k@�N�Cj��)m�m#�{��w��V�q�(w��)�3ԉ����G��l@ѭ2��ů�0�@i�����
��ʧ�.��!ݓ򸰅�<������.9%!��k����Ga|иQr,|���z*d�j�әj"!�Id9Y����j��܌��e2�PN����	lQ�.[:ԫ�_RX�R:���D�yS���2�N��C�&���%�!�n�6�>�}o��FiK�-+�A��]`2���=pdE��5�����)��2z��HJf�;�J閪��.���/���t�O�H�b��9��BE�G��������L4����]�}�W�$uldU0�?��z���s��������J
�َ42w_�K����*��#K��W���u�{�V���t��o5m�����r~o��00	�p���g�ɤ�� �ypn�L�/��R2[s�'m/��Ǒ����f\-���>Dp�-��R��.b�>����uc+�PѴ�1dܙ\6��k'��^�O�Y2�V�gT��Ǒ�6��z�]Z�7���\&/`܄��H�I��m�]*��������1YNzMl��s����6V��~�:5;�\�����q3��A2���;��/��̰#У1I P��(�[��?����b�Hçc�dUs���n�:,�㟎.]>UqK�t+�$���Ё'��E2
3k!']�~��u�gz��������k;�cg�㧩����UҞ[��[��\S�]�p�[�<�����杠�W�b%	#�	������pN���	\�4z|I��~�ْ���f6�$j���Ƹ|T����:9�]���c^b�w?�t�O�,��@�����/ɝ�uC�}N��O��&2��Ժ�8F�G�Ȝf
�^r
m����aD��'�Xq�+������ΰ���� h���Ǽ)�n���X\�{��@�?6���+��<��c25}��^�a	!zR���^����F�B��BNnв�~����������K1?kا/\7>@pN(��ĵs�����Y\�n��_DaA�]Rኹ}�	�<�YidT3��)�9i.�ȇ��1R!焹A�`%�lNN��
�p��@eÐ��:�b�N�K�v��#�����#�^��>��I��ɭ�Z�$ZR�<�2n݋�����T�dC�������$TA�,)eu��dv��|�jX=1K�73��J��1?�B��qC]Z�sh�`�33e�j,Vcu)͘�ei\�N�]���W��o}��C��d�Ii��{�[���C��x�A����|d�Ncj�u����	M�1��W�%��d�������a�����<!��i�F�Ⱦс�ʤ�d�����q�T���q�Ob�1�^�5i3w	��Fg�t��
M�����d�������B���"<Ѷ	�;5S=����������0�۹	��{q)�x�g���]=(޽����>� ҵ/r�aD���0m�'R+�wy��m7�>;�ۉcƁ���p��6&R4և�kk_��s�����a���1w@Qz�,q�!������<Ϲ��>"��T�`���(1�!̒�H���>,��y��4?$�ƽ�FR˛:�r؍2�t�>�:�]�.'x�:�F���sch��xYJ�������\� ��1��Nx%�f��*��%�P��Z�П��Uμx-g�����m�a�
S�L@c�;��P�-2[Y�l��P�����D��#�	��]�������H��+��F[Z��W���p2����G���=2���u�v���q��cx��M$	�%aT�z�ǵte���Ɩ	{����/(B��:_(�Ú����3�\$���Of(�#�\���/;P[�-U���ނ���n|�f�+;!�
�#��-���	��g���X,��E�� 7��ҙ���0UV�C��H��W
Qn�D%�_$d=Z�*/��<�̽�BqpC0��@C���׿��}D"�+gNH�Rʊ���a�;�'[�����������//׾� ۼT�Lk���G�Mfd��٫�D���B�Nx{��T.����JUc,�7�*;�����J��9��y���l�;�6��2!�(�^I����ņ�v?U~7��㙙�Z�V3W�k��o�ȹӧ��^#1�"�<�?\a��>æ��� ��U�	�P(�����{�aQzϱ�q�pV?�o���$\��e:���Q;��iA��0Ҷ-L��E�
	�?k�d�uk����l������f�,��ef��v�%n��i�Dbn�`�G ޹{V����/^2#:��0Hq��$�I	�� [9d�R�ʀ�e#��o��v�A�x:a���M��i��Y{�jY	)0�R-�W�����Z��ętr\��D �~����A���F�d����̍��� υaｏ[�F�ҷ���}���p�r'x,��q��^ꮊ���������Ma70�`���}�8��	:A�$��V��y�>��lWj9��䟌Z�p��PI9��_��#�$���cb�1&��s(��,��� ��]ךX�$�|��l!�� ��U0�,u��ƚK7�a(�ͪ��iO\IjH�]��z�C
�1���3p�JsN�qf�<��E����D��v̄G��Q��#��?�L��Z`6{�ZJ���D�̫����QOz{�u�� ����w:����y��&��Gi�]OT������l�h,��^��cǫ5�ݱ%V.�I�5��ɳ$��Lx�1�N(����N  p���"i����s��&�i/�(vu�����c����灴/4z��=F��Ԯ�1:b���������q����d�Pσ>_��N$8x����pg�x�����b
�tgޅ�ִ�8�ck�R��Y����{$}ؓ�\���%�L��fS����$�Ql"M��_�j���^��ik���}��Q��Ĩ�~��8T�?��a�
��6��'J�/L���=X��s���oQ�����I�õ��2��~��'h�;Kn��0f����LU^S��F9g#�Y�J	�$�
��o0K��v��W���?fp���񧧖�"�~�����6տ�!�Nl4R�Wc�i,BF��J�#2�i�<�f'�2X�t9o����ܿ�Vr_��+�ׇ�]�6���|������^�D�73Q�6�]u�'�����Sa*�O=�;Ҍ�hӊ��'��Ǌ���l���E���N��'ֳ�?�P���b�r�x���<����?F񼶋�P��F f����(5��f�~Z</l��%�~t؏�=LVpJ��_أ�(4���
�'`�k����W��.H��󽍊p�ey��ҕ��G�0�2gl������3I%��fN�=eQ]����;�P��� ��W㏃����&`��t��Ҭ���{2��!&1�6�C=���Q��M���b������\��?�|�1�ch7D<+��#XI�N
ժ���OY>��$3��5��{q���Ƨ�?�Fy=��Â$�>��LFtФٽdI�9�G�h�zŦ&K���P����@/�{q�;
~T��J���럅p7��E5b��)Ak�,(S��*�3�@�N�·��#���1�[��W�)��L'�_R�z���(�����:.�q����4��e�9Y��双��4ZH��]�s
�DNR>�<R��GT�Z�n�y����v/I9������!�~��{��q��T>wE�[��"��i�ˀw�|��O���*�����3Ξ�nV�c��1`fp�o���zu�d6�@�2w��,7tS��o�#JO�����JA �T~#C��}F�
&��xӼ�f���๣�x�p�,����.���%��O/���������}g7�0z)l���V����@�W����5��@�L<�@ "Γ�4��<�wVU7:�����1����v�N4E6��6�=,#ϋ���-X��*���y?����?��8=Ͱ`A*:�.wtc#�@:N/A�3�:��ך�l�됒F�Lv��Ką�7����M�9��w�}��*�����F�9��@��y�#s��|�a 5�/���={	�7���}�O.���H�]�IA�?r�{r<'F����+������+5�&�0~屻�9Ͱ����q����́�U+�(��3]첌�#̏0�H{���iI#��l����#�KZI��>Z���6����VaK5�j<�3��\��JC���y�h�-~S�׃���13�\�na��gĘ���GI0��<��ޘi����`s����G'e�	a��BX�2��xp�Q�Vb��/d5� �%� �5�X�<��]Oea�C���0�YKA4A�Qk���´{?�mn�L�`�zQ�em��Y�-�ʹ2Z�P%Rj�E���Z�7	a?N�ӛ��k��R�����}Ok�9`59�M�:�wK���z|�&�ZթF�)EP����k�{V5��Q��P�m�2)����fy�А1�T��(�'�&;w���!����/�}D�n��q�jY����&��?�6�5ڎۤ�=��7���������h,�j�zYqH��ն�m&K�۷{`�]�];���s�NA�m��O��Ф��v,��\���~)%^��G^��Wv�:�8!v���7`x9�Х�_nߍ��i���c�w�,m3��ce˃5��0^,R~ݍ�0ɌLv��nȽ��5�si�|��/�Y�.�
F<u%���_��O���^B��p9�z�O=���f&�*��搬��ߟoM!�hk�����NH�������>�VM�����9������m|�����V�.�|�썯f�=�Z�Q�H~2��%C�ɵm�7_���Q��E��&�|wC�[w��x3��78��NeV�o��UT<����y�� F���(o��}���Y�� ����G���yϥl6F�&����[���~�}�����)��4��ɲݦ�܀�������y���-�(䛞U�6�A[9��,�_��ѹat�����Ć���~���&#:_��5��ו����~���|O�O#3WJ��'��Ǥ�~���������z��M��^�� J�C㧷"'DXn�͙����D�⃘�`c�|[t�鮢����W��vqF4ks�N�xp�4 �v^6�x�4P8��R�	Ğ�d
��<� �㾌�~Э��N��J�˚�������߆;�������)���ۥ�3*I���f��D1���~SHB���m�����rW��f9I���^�E�ٺI��L*�-1͹����h?	&�j�����p������U�K��Nx�o�Hc\u"e�+�Q8���bՌ����WbA]J�T[bl��؝��V��Cc�8��i�Jb��e���D��ө9�Vrѯ.��N3X{�{���5C��Hu<g!�ځ;,���n�_yՔ_�|ٺ%K����ݝ�D`�Zpj�"�d�3Ĳ�Q����}�K��z�
�d��@>�x(���/]_�3kf�M�Yʿ�'�v,Ֆ�0n���fA|'�m'!7o֬���"�	��Ce����q���Wt݃��D6�ZT<��P���ƺJڈ�:I;ѿ$$���	�Z0HƜg#�h@z�ê�9u>yX����݃�X���ĉ��z����i��?}h�����%���!�?����n}�L��em�6���9*�[�h�r2�.ES�e��i�������������àu)H���{�{bN��J�{���I�W�ڄ�Ԛ=�W0�V���2#�9^��5j���ՎbWl�^̡p��;_�F�.ݽ�C�Wg�������<�"��6�W7��7mf`�4�����+/#p��N�Ws��;�����C7��F*ޓB!�{�{+�Q ��U�s��}�zԌ�d�nE'��Up+z,�8|,9�����~'��j �υ��ߨ+šѺO8��㏕!j��H��y��Da�I��ղ4�O�ⰷJU�6?���YC]�*��rm�P�դZ���-�8mA���9����Q�����N�,�����M��)�,1J����枘����ж�;Y<A�p�>�d��kñr���X%9�X#�9�:�� ��Y�����A�l�V=-�1�Lu9#����j�̜�Ҥ�	I�Z�E&>���2қ��g W��	��E����`(�7�����ǂԂ���2
ء!` �������Rg��X��Apaj���,�3t�Ugi�(�%0����b�L�����lXB2�{�E�F���V@���Ʃ���s�~9^v���ge��n����GF3X,�x�EW`!�qpq�a�_e&3y��`�a�9K<G9�O��\[�O��aq�jwQ�)t���''���\�����ҳݒ1��K����2�t��7�soIݵ<��q����f0n��DU?;�;`1Ʀ
��g6D�_#)fCX�31+�HHژ�r$sOb�ѻ�����m��M��Ν;�O,�<~�Ġ���	���<5�,��M/G+�0���x\~�Y8f�z\w�'��El���o��.�@¶߾�N�x�͈<_�Lz�׬�/]y���-v�����0���H(>l����g���߾K��{���Uo��~���}�������f���fg���g8b�4�t���ވ�}�.lX�
�����7�J��8���YZ��G�YY)��v�}�9ߺ�Hl\�F8�KԘ�ל�F�ĺ�	��z�3:%�W����sx��'�<z0Щ��3��سg�<��b�K	�?��3��O��r�/lj�|�w>���~�<x��_�>uí8ԏa��F���SO�����k�N\����ݹC�x��1|>�v�ǿ�8����g��Y���o����:x���?�^����]�ƞ�v���x��'������~��n�ޔ�/s}��'�+���|�2���G��+O���	�^=�����{��U�i��9gzӨK�,ɽ�ml�������M���@BB�	l�lI�}7��f� B�&@��fc�1ƽ7Y��FҌ���޽�3b������y����ɚ3g~����]�Q�%�|^H�:-�#��!�Z��iHY��|S�To���y_��kV���Ϡ�|���-��*���d�t�}������P5r����o�p'��Fp��&,�8n��;��"X�V�Y^f����
+�sE���kم�l_Y��D�Xli"L�r�wz��Lf���z&����.Z����ǘ��K:ގ�_�(֝��qB'��!ӌza�NW��Y��f��� �����RZ�#����t�N&+LZNq�^��lIt������IC�t�%jE{L�Z:9�he�fN��o�*������=�����ɡ"r�:�]q%��Sd����i^X�Y�. w钠":\�ԄeoN�2�a��FK��:�"�5R��ENm����w	�T����MB5���J�0�a<8��NL���5h���Lc�v	k��������xRsKt��O�������{o����'��cu�4z��.����*q����+��Ϲqr��f*Z�!Δ�r)T�,x�,�ZC�Q��᪋a��&<����`�^Y���}��b�E����x�g��<,��?^�E�F,9"ĸhu�X�V�F0v�X̘yrE���������CRЙ�r�5W���A������o��=,r�"���/?�)jk��=���}ｽ3�L�?����6���y`A�&G�=����i�����t2�\6�sfMGu�BV��� �UB����E����<�9�`�G����G�p�t���P�ů�%nj���p:��To�؃'NI�������{'�,�@��ϼ�
�{���%�nU	%��$<��9�g��w�.��M���CG� Mݿ�1��n�����D���o��;�އ�H�eᒕ��߽����ؾu��%�[Z�Ʈݻ�Υ��g��\[�*]�ȽG�1j�$�i��1�|��N����כ"��톷���
���� �PTP0�r��T�u՜so���V�?����S?�8[�?�E}ʆ�=���X�\R��)�CX��J�"zu����q��Z���X%��PM^�[��|� �N�=�8�b��s����#�)ƜN�8��y�Q��BN��1���;��P��0�����r�7�d�H���c���D
W��7�n����vyd���uK�]fMU�tU�QTUE��=tQ70f���Ǣ�~�t�������Q��#�lS���5|&�'�d��ԩ��#􈎙u0���q�uW!f��r ?��	�g�j�<�|���gYp�RN!���$�kw��r�A�<�č�+^��~9�~��h�D�%j���f>�l"&�,<��ŝ<Cp���~��"�����`�d��ak>�tہ�i��@�W�����w��T�Ġg�oVY��Y����a��6�����4ԁ� �x��H���C1Є��3�D�,9�QH'PC���BPI!ֶ�ZW���&���?�'�i��q���+q麵B�ڲy3�}�iq:T��(J���YsQ�F,�����6�Cs+���ro���c$]��������������
���/Ha�`�~����F��Ef5�������:�#Cq��g��ޝ`�����]����:�t���K2>,�+��h�c���=R�9%s-u��%0��� 8\8)���9�o�-{�[�)w�� �:���nq���#���q�4lH�FN���e�N��#�Ƣ������e���K��0�k�\xf����}-�P�������]*|�d2!k��σH�B^Kmu56���=�b�h�	�b��k��o߆ζ<��C��D�QUE{{���3��4�4�5��5� �ʨ �p�{�R=D������\���Nq6��T�MY�7�J�|A����P�Q�_pyLmjxkż����k֞��Ϡ�|���-��*�N���?l?zo��Y�!��zK�+fs�`�;���|n�kn���j4����j-[:k��2f	�D�P�����C�ЗH	���s�Q�bV�D�����i�a���X]���@	�]@T��5+q��%�z�d��;����=���^x4�O�(����.��oF�����F`a~ȃ��n&��������U~��yg���ƬY�����DNC�s (����fxCQĒi<vB$n���g'�WUY���zTE�bG�`���$�Qw?�h�P�/p�go������޴����>�ߝÂu�D���`�)r�%?������g���G�y�Rg�t��e�EX�4P�fQH��m5���V�iN2>�tb n�&8E(�gWM�huʹ8���rdCb��0z�kP=$s%���D�$5:���Jhޠ���`@K6JYG+h*3k����.���^�4�D?����G���y�V֣�e:*Z��Q�5dţ�+�*�ETX�(��'Ӌ�/�Mc���G��]�v	����E˗aݚ���<���F<������(�E��Be��f�Ask�e�~�������e(>"�ѓ'��;E�84��U�_�/}�&�����6���,����ʛǎ����;L?�����7���>�u���������1S-���2bB3D6�r���TUTI����$뜒��B����]Hm,^2��%N��ӝ07�c���� ݽ����vV
tZ�a��"Q(b UĖ�w�`['t�����C
��;��E��*�ٗ6���^�P.C����V�D����p.[��7OX���r�<*�kO$q�T;^xe��P,��nw[>u�5���[����V��&�c�0H���� �9�N#?Ǽ���]��G��@�1H*s~�Gr>�O�@F���s%�**`�*`��h�r�k�h��{}��Ew�ݡ�A���O=[�?���JM���'�����T
�jd�}��K�g�#㶐AX/b|ԏ�c�x�4z�@�񅉬i�?����m�{������-�h�!��~B?hN3b���Ch���%�=�9���HX��Un_��J,��"K��!<��O�����L�D[�z��?w&r�aѲ����j9A!���fRq�vu">4 ����K��}��ޔ��NP^�Lw�S�AT�/�����}�>�GPUY#�+���9Wv�-c+q���w��T����ر{v��/�h���?w:���PUFNxq~��;���z�� b�"�a�YϺ�ɂnG*G�!-e�nV|����ď�ϸM:��ؤi5Ṭ��l�|^:s��g���F��Lhvn3��WCe��]�y��r7L��׉ML8u��,r�o����ny`��P���M���p�=I!_U7�G��钊\I!�	��r	��i��Bƣ婧���1���a)^�ťO؛��j�P�) j�P�C�Ƶ�\���F<�أؽs��a���X�p!���غy6<��X���_	���'N��hU�܏�r�O!���UȽ��݅;w���#�rzk׬��?�iT��������}�"����6\0w.����=��/����F\�n�0�����@�J"7�֜rB��x=�*k����rK�x��4��*����u>A��,F�>�L�h���X� G䪿?&��ށ~q�㪪�ik��&�"Y��O����p�T'2Y]d��zfA_�`>txꅗ��/!�+���4k����^(߆fC$F6VWaά�Ҡ�9�]�rG�F��v큩�DV��}1������m�����ىcGc0F�?0D�ANd2H�����I�M]c����׏�2���0<?�44�#*:Q1�?3�����
'�M�[/��a���-��wnX��38~�>�c\���c\�ѧ<ؗ\p��Ï���)yƑ���`f�b#�g4(uV���O�����eB�Q]q� F2C�4:9I��s2��A�]'�x:�I�"�<xLǞ��LN��vl 5I�j�z1&����$ƅ]H'�8x�(zf�a���Q�,_�5+�BQ�7�AHX������9�be'�Ab�#�!�Mr����,���THΨ�S�|a����EK�p����O�76,.pt��7g.�/Y�1uaT�m�+�c�y}�Vlݶ]N'����s8���(i��Ǔ��珠e�j��Z&�(�8�;0�p�l�eF�ݬ�;Mg���P���T!��A��!�PB1�Afd�)�7Qu�z.+���v%�ȑyP�$��q�#����J���g�L�p�{�tS&�ݭ�I3�E�P`�ғ��z�FQU7VH�����/�\!�*�.[�W1PȦQ�D���
V����x�/0Z��.=��_CT͢�D��H���W����>����'�;�ĥ�^���_��h�m}�>��8��\���{�Xܲx�%���������j�,⇎�}2�E��ǪUk��}�h�����_��		�|���V,9ܪ�=۷����H,�	��0e�DL�:E8D[�Mϴ::�ь&N�c����PQY-�^�:��A�0�i5L�Ks;���X�3����0M)�,`D��پ}���ѭ���J�SN躢a ��ɞ!:ى��AIX�D������?Y����~?�'���7e�%7�_��S�,�Xz!̝�Gy]=��A����5�p�Wa��C����pY\���W_���N��yv��M
��Ѐ�)C�1�>yʱr-�`���W^�����+�u�wleG�8��Ş?3�#&@2{��Ί	M BѦ>=
��G�<�_\�xv�l��w�;��f��}ָ����j�!"6�)��S���>zZ����O~���n��v���*|�m~����������������^�7Ϫ��˥�Jb��r�Y~�sE�å(N���誡j.�NQ�MRU�4-�_S�E��66���2�!�����.�}����n;�`�;8�@�%I8�$r�!�=~��~!y4�!���䴕Bi`�O�    IDATnBn��!�6�,��4j?��D
cU���i�L�"Ra����p�������!�s��.��c�q����ĺ��a깍�I0-�S.[�W]�^��ښJ�'<�xNa��=�P�@o�L晑a�S	�q�L[R�>�������&�=��؉��*r��L�HG�i9�j��`�ܹX��<DB"�Fwg��S�#g`���xs�V)PD)l=��\�/��9)���=��cf!�D00R�)tɗ�q�]��:+';܉�UH�#�*Ip2�pR4a��H,���{�g���m�S
�����y��n	ވ=�]��0���|_���A�tg/N��B�PR�8��"U�pE��6�[݂D����m�2�uc00�>E^����8�F^�Iң�hV<yg���� Ǧ}/��:43�J5�pi ��qx�n�j�L�>� �>�x�k*֮]��W�R��۷�'����n!��ܙ3����!�+Z��pR�@�4�<�[�����ڍD&#�ʵ���+7�"<����2�'����n��.��F:��/<�ꫣ�p�"L�<	�Ԉ��b*�u���Z��E��	��j��C>�BE$��alE*�[�de \1p\��'*&����;���$�7�|G�F?a}�>�Gh5�3�,��{�u��~����-�{�X-�c^� ~ON�����ψV��҅q��_�����_���C��2����_��O���>&k����Iⳟ��x�mx��mx��W���.����&��p��!'�<��N�I�|/�H��bd�K�}������_����?����#	Y���G$����c�*�a=N`�mf�#��")J�P<�e7��:V��U�v1ƶ�0) �
�r'������.��R�R�kd&2�RM��ض�3u�oۦ϶,1T�=�/-�E�#�ضB�'���i�b+�7䱫hrt��!��2.b��ؖ�33bZV�JB��4id�g�n�4��@e�g�ԣٶM�k�H~ar���ʪ�_�|՛ʨn�jӇ��_�5�����w�.�o���<�	y͍R.�tWl�k=�\�����{@�WE1�Ɯ�TAEA����Rѐ�U�KOvN�sy���s�aA�t�����9Ne�D�Ew������c��r�\�r!�\@O� �~n�젻���ft�W]�O^{%<�%?�Z��p"��RI�@�{K'���8�\*%�6~�I?sb3�5´g:T�4�u�t�t���K���q�&�sY?�&N��Y�P�(�����Ϫ"!1���ڛ�M�M.-����u��I�Ł�>�Io-�v%���N/Y2�iӄ�(�3[^��b�ϱYٚDf�e:4�eA�Q�g�I�PHA522��Q�_+�.���
��f�>����-Ho�@@��Lc�a��p�x::{Dڕ/�r��!��j��c;���"l_�0�'L��hM�=#��2e�r��zA������*����/5�:�#�������t��mfQ��������b�h�YЏ:T6T���K.��K�ja�]x��a�.ULe8I�۝�� _��w�%ާ�������C�HrX�e���/IA?r�$~�?���aY�pu�~��x�5h��F�߇-ol�O���2a<V]�\��b��B�+%��z�싄`���67cض0\b=��X[���_�z��DX�ɒ�o�
��@>�@�S@M�D������=�f�k$�V���"����X[��������w'/^�T.�?<�8�x�%1.r3���Ur��S��|�L�Њ���_a˖�dUG�C�&O��������ڀ{|>�G�z�MIA��۷c��;��?���Ml�'�6K��hA��6`�f�I��gY��Phnnƴi�俖�)�\ѕ'^Aϲ��;�0��Kh/�A6@l�)�$����&�ֶL䳭�KE��Ȱ���~(�OS��(M�(�es�c�4�CjӤ6��DI��
�wHŶmL)����߻�����S?�ǚ�8#���@g�����ɼ�j�_K��S��2��`�]N��|����y��
�R�d����,^��<�����	�.��{c=��?���s�1�e�;��ѥ�^Oj���ƈH�/u��,�L^��Rr0wKZ�n��Ձjɸf9�@�(�6���i˟�	I��7���5+�r�D�&���s�8���7�\n|��u������ؒY-w7Me��l-s��{:ň$�A.3���A1fa!��:'@��9���J{uU�͞��l	}�:b)�k�FW<���C��	&OC��f'����,栔2���{����[b��ж����'�{w�!�w
���o"��$�HU�ʀ�5'�Ҕ�kѰ	��KN�^锲Q�L#��_�|I|��^,
�<���O"���J�E�\E4�<SBu�#�{�ӹ�����G��P��O���޽����+f5��uV+��0�b�;u.����pQ��	��"����T*�\��b�M�O���4E"\��%Aq�H1�t8��iP�����it�6� ��>���q����d�+�x���q`���I���˱|�Eb����x���Pb��W��N��E}�
���#A9��@�_������<~t�FGo��^�_��b�k�^����M�|^����Z\�x֯Z!.ov�����P[Ō)�
���1��E4��5oh�[����j$m�bI�|��0�T��0�B�h%��)8�a��N7@�����uؼy3�;&�S6)�zǯ�+y�jq�k��y\�����ez}��������� � Ò�GC$3�L����^���?ñcGPQE�Δ����_s�~�e����;�����!��>���o݁�{>���AG�I�Y4��bxx�O�;� ����A"�W<y���ɓ'K��i�D��L���9�g&8�3���q ���Uz�]/�4��~�Z&�9_��I��W��Sty��*�������0�r��� ɯ���k%ʁ���p!�Y,[A��#_q�F� ����/8���K���A����Jb���ճ�_9#�Љ���ICt���ߋJC7�+�Juuu�\ż�W��<����ق~����l;�@���cw�ˠ�ف�@?|�0���h��E�զ��Q7�IH��Q}�iA*^�Mc;0稳�]�7gA��V���;P*R�ŉ_rVS}%�Y�
���0�������ǻ��a,��!�q���q�� ��G������g3)t��Ʉ�4�B6���^�ӽy=�y��h�7���f:�H��_(iq����'���m��P��&4M�*:^��y8eFP�,�V�p��~���k�VѲ8o�$��w�XC_��#��N���-jU����9���g�p\\�6Âfڰ����D�����C������̍�m�l�����D\%4��W_�ƚ��GN�af��$�51�I��� v�ڃ��~��fښJ�l&�y�4LĲ+nD�Ĺ8�9����K[�Z.��Ǝm��l86�\&+�0.��rj�m��]|�P���CL%�CD���U|h�㷳�1�b'B
׬_���*��p��iNX\,X�u����ְc�{x{��%�	��$I���eŴ��E���ũxpH�N��Q5&N��@8��'��
P?�	�]q���s�^���5$�<�w���~U�d��XD����"dFޗ�>�qY}��p~����?X>J\eq�XU�A�%_@�{s�F�,JV�%e�cqW�f٭���;Sg1��&�t�(�5�Opt�4\�Tj��l����IKA�?�@�O=�'<��ϲC��=3�m$�ru��2_�鋈����bϞ]�Q 2�󥦱���w1q�d<��+����II�v�W��;������{ݧ;�~����ޮn9Kx���;zt�鐯���,���;�<)�3gΔ�{�|��Q`���Bow�!A��PJ7��z�Xѩ�?'SK��T��+��G�S(�3�~�?a��rBʫ��d8#d,K9�/�>Z|�Ў�5}��?Z�G��I+�ܣ͆c�����kykW�˿1:(�^�N�-�l�Cuu�?�xݕ�Uf#�u�������e��{�>�ے�b>��e8E[lT�*)B$�xH��	ML��<IX�	)��N�'���t����9����#��9]BFʓ4w�d�MѠ�Ua\�z9�/����:Ԏ?��8�vR��׏��W_��]y)BAgGFs�<}H���4�4:N�@6Im�c�2�G����.�h�Bݑdҙ��i�!6��-E"�c�qtg�ľ�$t��z�:�|��Qt�Ǡ�xTQ/��h����l}�m��$G(|�9Sp�w� ��}��z�����1�Qa��3m�΂a����?gK��Z�"n���
�L�l+�-�3#��	Z���+3��8����ڐ[lO[��KCP�P/{�hE�L����;O���6�ܹSX��&	��u�.M�}g-X���~#�����Ɓ�8oE�QUS/����^Y�p-�Y�nɣv��z��L�
dKh�������#Ì�C Y�K�(�N b���W��	��{�ǎɮ�&$uuu�2q�|�C��"���//�$I&���H��\�h�S)�$��th��qط�����'Oy޾#���1Y�� �45���OV�K�%:w���
p��sq�%k0n\�H���aly�M�8tL����$5OC^/I����Hg
N���<74�s9�d����Ti���:1�l�~��M�󹌳kW��o�C!��6�KS��L.���OfD���%ɭ2��_��'�����_�Sz�#I!�It�i9�����i,���J,:�<��8�ή���ux|!�����`!�~}�����vQ�p־l�J���;����x핗p��$|>����8Nwtȵ%��Q�rC��1��4��
L�0��������ڊ3f|�r%{ʴ�Q�4�N���cIJ��*�v����%��Rn�X�e�X��G�/���T;z\tBv
7���\���]��_~�	Y���:S����#$��G�=:@�)���Y�N����韟/񛐞�Ӹ�B�3��� �]>O���^2�|�T��Pw��������}%���Գ��ޯ:�W<����!W�)ǂ�NC�逕!$Z�����^v��,��.�P�V�RQ�Y�'�>����s� ,2�� J4C���F�����Jٖ�=$Z��g�J�eTq(#쩙y�T��~�ܸv)B*��c�=���vҳ8�1V����S�_�H�C�c�LH�]7?؄�(���f�e
����Y�HX�ϓL�8p#!}uu�h�4CYG{�+��u���1��pE�0n�t���b0�mK�_)��:�J����
��HQFR��]<�q�W�99=���~��y��Л�`�*�9�t�`+�kf/L(�$'��5�OZ�r�Z%��RPHg��@Ԅ�/������.j)�b�ji����֩@˘��6�e�T4�oE��(�ߌ3-$#سk�n�*P��+����`��w����Ϣf�d�|��w����w�3i"o�����3�в�	j�}nI���5cZ�-����a����0�MN`�g�N]GP����FNKA_�|�L�ԡ�vw;:e۔C"a���l��Ģ2���I���ǝ��
#�ȑ#覿Ak+��J��x����	��2c�Ȭں���3��:|��]`A��k�;/�"��>V��W_u)&Mh�5L<6�����{D�x���.�F��V�IeE�悃p�u�t��m���ɓ�y~k���\������e�p�왨G5N�^�p$�>G#���R�Xhy�3D��s]��C7���
47�
��?0������_�P&�咩���/���~�8nn��z���WA��l^X���0�~����fY���B��`ι��7��#������KP�h8$Ll�O�A8N����Y�)aljj�ezMpBw\$Gu�IP��������r�w�c'1�A��@:�"æ�d������|�T�g�c;��9i�-����6˰��`�|�U9ٗضe��Ə��ùmw�s�˜�)��=��RT�qp~/��9�sMO�;�B�#���zsU"��i�\�[��h��UQEQ��)٪�����f�4���j����+�V�-3k�vFQ�MՎ�m�p�������|�-�gp�~q����v��w�S �lݓǡK(
cŇPU�Lؔڠ�E��O&��Zq��5 )x�����6 g�7�.�p���WDd�*�A'x�9�[�z��;d~�H���lTE��?sn��j���<^ߴϼ�'���4PK����?���ť���;�����P1w�m'0<�+���� ���T�C��¸+���0�B}�X�4�` U@oZGwJ��ǻp�t)�OU�Սp��r@�UE�H6�6w1���w��wߓI���QV+���/��E�����_��&.X���$�}
y�N���E�߅�l*��<�)���D����	�C�z)/��!��
P�d���UL �6�,)���B�:�\L�>���K#���yOW����ߏt2��,CLJ8AVTFp�����/���0Tp�+m�=����'t���G!�ICO��.8]�௭C�䩈�������5�9l�ZEy���R
z�� ��)��8�X��CR��G�m�ӑ�)�e	i�
�{��j0	I+��)S��h���yc���oű�m8z���ol~L�]��p���gr�@�5�S$(�u���8��=��o�?n/Z��.��i�����q�A��ݜ��=7s�����*�O�%r6N�=�xj��x��WQ���㕢�1��vI�77~+W��_F]�r.6���X�]������b#��ĐH!��G$�j���B��'�ņ�oIY�^�mG��&D"dA����ԉP[�Ͻ+T)��O���;�G�RP$�4_���K.ĝ�~￻o��g��{ER�P6~�=]r���2�:i�PCP���'s��X��ܱ��������k�D��]�܇�6�Y���fJc��s�r����r��n��"��
9��rY.��$�A�R�TW*r�����۔��\!�eJy����|���jyhZ
�]d�����2�7�j�*���+䙒�N������JAQ�Ǚ���(�F7H��C1UM�U��䲔\｢�����ۥ�*
�=�bۺ�cX��[~����uK��V�T��P�2�8k֬rf������-�gpv��Gv��݈;�@���'�*0�a0��,��4jT�bk���uk/����-{�����3�^I����? ]7���"yE�C��ss�r���b�`�yЋ����'�ǹc#(�ǎ�����|p��c���x!��Q__-ӫ8?QϬnB�B��GۑC�F��X_7�ٔ@N� =:�-898�I��@�Â>�1$A�'�c��n�>Ս|�Fk_�@��b!Z� �Q�blU�n݌�^~Mt*�ˋP8,��Wʤ��]��7���Ϡ}DR�byQ,�ݎ��S�mF���f�#EB�:�\z:	�S����'�g� Wt��k�8R}'�Wr���{ %R���kK����2a<f�:G?Nq���:,���!�ZFjX�\>/�.�H��)}"�+����A�θ�_
`Ў�m ��N�\��H�%5.�_��ʆzē#�'G`�e�h�!	�9��D�e";�����L�#�ep��s��������^;$LJ-�)��o��Ж�S�oI��%LKW�Q�;�����'�v�4B�j��w0����7svȴ��p{c9��b�_ ���
�����
��W�^���cdB$��?+��}!c���ZT��y��2��><��l�����eOd�(���=��u�bŊB���'z��bk,d8�_��T��|��O:cI���Rl�II��9LWw/y�9�?��D�M%�"+4%;�����V�Z�L^;_��?4Ml��4m'NuwC�VIF9:'��˖�k_�	[�|�����z0��ɑ8N�>-
�����|n��%�ٶ�l����D��Yܥ�){+0S����a    IDAT�H"��Ј4-�n.�ߖ�<ׇ<lF{��H�/��P p*Rzy��	�7+^oN��E��4m�+j��E#@��U)s��*2"�TL��ִ����y�4m�[�<���(F��t��-��T��Ƣ��a4ɯŢ���G�P�ߟ�N�X�ܱ�,?��H�Π���Գ�.��<~���v��C��g:z��V&/D_(4,�M*��$�`����aͅs$��{��c �AF���qbH�K��N����+�S���#wU.qEz54FC����Xw�T�����G����&�n�mc��X�|9���厐����TzD`NZ�=�����)�<�8����a%IU�*i�B�����2Z�	Sg"gi�Π'UľS��}��;�H�`�5� �U!q?��S��/��'�{�Ǐ��`�E���$���1���'^�[;��O�7��@�ˠ/�!a/�lUi�Zd�#󉇻��^��k��
y�tI�3K���J�����p�aԄ�Pj̽<'x�:\.9���\~�40���F�����>'T�MPG�v����O��Z��M%Q�5t��}'q*n¨h�Q9'b9�7r%rԝ�B���Kw3Mȗ��JJ��/:��B���W5%�FA
0�b�b�� w�š6�G-\��\!em��z�;���9(S�8)�L�����0PV����.\�X��h1:
�����ʦ7�Xd����2�\ԏ�G�|�$
|?�)�4Sb1��dq!�b*AP�(i`��ɺ�6}�H�$�@�a*$Q�`�!*��ȑ�F��m	<��׋ �����T�N��?3�M��l�ĜHU���LG�����2	�	U2�K���)lޢ!�⃂�1�����8t�E���C����T>j����;�~�*|�kQ�{`2���_h����ko�ݻp��&w�<�Y�\����-�˖����Y���#�=����C&t�%d��v�3,�|M,ޔ����?��F��"ɤ�{���E��+K�z�$I���^6IT�D@�S|3�n�UG�O�<�7�.�p�+V��|���W�lA?�[�_Ot^����aA/X
�t��J	:�A�ξ �-y!���<",��<�_p.]v��o۶�<�$���L�[�т.$�t��&�#�|�a������^�J4&�Y:|��J��gN�g��c#��bρ����I�U>EÒ��n��rp�����]3̀����[N�8&�*�}��v	l'{3U�hNQb���%�� Y�6�� f�slo�=��J�xW?�;������31��E�Ei�:gR#�n9���&l�����W�*ڨmj��|�sX�t�h���8�_?�Nf\���Z$�
�a��#_ɨ�4�i�D]��r�:�E6;��E�8���*d�R��5#2Rй;��@m���g����#o�{���Bɏ'y�h���	��A�9�	���n��.\,�(�U�9r�nG79o��f�#]()	����ʝ$m`�?n�vv޴e�I�R��g���B 
,[G��ÕbA?�1U
�?[|^|�1"!�]Xܜ69�S�Q̋+Y��I��N�;��kW�СC2�������uؼe+,ՅYs�c��h�8�>� �R,|l��.a��g�`Q��F�z�@�:F�q��I� )����;%}>Ņh(,���a����>d��m�y��ׇ������Le��29��-�Ow�	�Mu�������G�@�N1���D]4*M��|��4Z]����(���>��������Di�b$�4\o���9�;{&�ϙ��Q̑���'O��ٳgKQu��x�/�!�L����e�l����;��{o�M�H`o���j�@��Wd�1�g�Rٲ��2_��ѦZ�m�C%�3j���g�fc��;��0��CE�W�R�rCJ��.ٽ`�컫p���X����>����+p�������]�<�K
zMބh?�]=0Sԡ+�ݨ���2��[Pt!`�`�0�i,�O�)�ȶ�v��c�d�BH�L�d�x�~��`���1�ӱ1��@�K�D^㶋�[%�D���5�cɜI�@:[�#�<�7_{�]s�2��x�C�	�0*�k �C1�uj���I!�����G�Z�W��������*��%��hh�4�@CL�J��O����B}�84�kFMu5�!f����QSS%����a<���xi�fX� .X�\��ڪ
��}��x�խH����ϣ;��w0C�m��S塨r�dc:���:�W�D��<)��3��(iT��h�j���0��ѓ@nF>�1іҦ��;���:'�aU�B�����Xt����x������ȉS�u�$��&��X`�Ltf��ϻ`{+$ ����t6#�~ʥ� {���1��#����ȋG�>gȄf���z`$N�*PĲ�*�3�<��ǎ|��.�R*zp���"�3i�ļ{j�iV�*8����u��}�I;�aԗg��Id�cs.�c۶m۶m۶m�8�m;9�s�ɉ�}ޭ�O�#��ꪞ����X�O�t�ѯ�^��������p��f)H�N����&�� |��U/4��sF�^�
š�9��.w�y�_��������cs����]?d�1ȉET��R�f��~"/��[��Qױ���h�_ܖ��!m�i_-ZA'�9<��+���;-�&/��Z��~�y%5�f5Q��^g���_L(�]��ve)�aU���ȅ��j0
��p66�N���&s���	�{ǔL���M�V�_��@�+�@B<#_�J�G�;;K1��3/^4��-��≫J��jec�b���`��� ���B'�yk {o�V0����0d��HSؖ���0�c����~�\�~��7����/��� ���?����Q��ðzK)������V$u9�����J�pV%T���X�j�r�d�1V�sF��&3�{���;�9�L,{U��H���ܺGU�I�����J�r���!3l���-���9�`;�q���@���[��ȱ3*Sq9��`)_�d�1��L��M�8����X�2G*�$�x��5�єZ���Z։u���#@Xw;�r���3�^����x�#�����̉��v��w5t�����a��۵�u�~H��}�vù��ڟ���l�E���x���*P�M�V:I�@YNex�[�d�V�2��0},a����$�
?��)3�I8����T&i�c�I�
k�Q��i*xM�4�Z4MJϽ�����O�l;����z���,����� �n�;�b�#1�8D88�����8e����U�e�Im����~ $4nөh{*8�~��n�|>p���Φ�wO+�G?},�Xg�p<I�(MY-���Dҡj
N��1�=��)�����lX�ÕƵX��<1��LQ!�2{~�3ba���ݠ���.�\��.3sZ��Sl��eE�8�mm�+�}�g�w�|�O�Qo�*��?G��_ð���?(3��#��g����1eD����+�����b7e	�,Y���]�Ӛ�'�_��K++�!7a�H� [�>�~���dy���
zsmjM��o~��x����o�<.g�]��;�Ҫ�H3剖� �m�^�ԫ��Jn:�ĉ�7l��*Á���n��	J�wj��	�WE�O�ֶ�X)a����L���[q@�xϻ�
���)1fY\ib	�	����0OU����ɸ��f����\^/b��aP������cبg�G�Ƿ�H!Ġ�%�ϒ�ǁ�������O��>�.%=~�wЫf\3����5 �C�٘z��k{�f0ۉ���[͟tx�q*�%�Ls���Ł~?�"�KJ1�E�M��H�{��]�����.�կ]w��j������v^6�b��'5:�.7��v8^n�(�M�R:Ǘ����E��PF�G#(����eT�*ˊ\��H�GlR�'��4�a�7��|cf��( �0�[E����#���z���:� ��v�<$�mH��G����+
y5R�l��_��6ݑD+0u lt��眽VW�$��i��kWxL$��11�)û6�s�!�"y����ˤ�X��Z��lj�V	&6�`��`�u@�1��p�=����Rd)���� RY��A֦�u��ơ$�n'��'�C�g�
�~:��C/�M�����VωE�4Q��p��Q�U.��H���0jձ5w##%�M.g��΍�#]��ndy�N%�RDԚ\_wT��btT(�C�q%���G��4i�{E\'�� 1�����UMCz����!��|���2^��ZNxos�p֩Xج���5�I��yT����҉�X1&�/���ꅢ�z`G�͸G��}��z�����q�X�+��Yv����q<���o�&�v����a��l�5
� ��kY��zX��~����:�׵Fh�l�,�W�4yA�Tn����y����U��f6��ф���ӫt*}��}�mwl���?�c�̞�o�ʨQ3�췩ѯ5��b�-��I�7�3���B~O�5� ���W�/I8D�<|�:?Yp�pZ%dhb�R!��)v(��ΏKۓ�w�i" �s�Г0׼/��,?R�0�� �B��SS��O��ϧ��*�;��ς�����0Cˮd�B�r�dU�,e؀Jĩ��T�A�(�R�-bQ�7� ��.�+m윸x��!��C��m��6ހe�s��f�3��j�k����ݦ�#�����8K��F4XkI�M!&{0��|VL:&���hh����$1�;:zH^��˹����P#i8
>o���l()vr˱�n��4�s��k��;i�.@TYMά&,=Ґ]�X�*�y^����$BCz}�Ox=\�D�f�.��:��F�c-�]Q��B|��'TPm'�1�����k��g���/י�
]�S���?R�r���\��!7~|P�睲
���&�\����l������eeĕ���8Tѱ?�4?�$8KF���2�B3Yq�z�����=��B)iÜA��,1[��X�Rx��������/}k?B]<p�tUT'������h_ �d"�ąe�
�}�0��V�(%u��K�e��'W����8e�Q	#.��jI��(JY+�i�E(ц��>����������)T;r	��0��d%��͵SH�B�A(/�H�t����W�E�2L!I�ݥ`>�e�9�D0=���5�t�i�U*Z_��1��b.Ȇg�,S�PԚ�*���cP`�r�H���o.1|��気�K���@�:]������� �H�v�_���n�5>�鴜
|���7�X�nzn��M� 
�+���qMÑ�>��:2�=�Lf�����>���h�ۂ��@+�7O=z�~ ��������4q���v��"�:-%T�c�g����Oa@T�FPc�tLi4�5�Ba��ދz��Ì�E8&yK�+�;#�|�{�E���(���/X$"~��^�{��}��;������Z�\ �����z��rL	�V���˘(TI\8��F���voX�.:���Hp���^lU�GK�pN��B>"� ~���/T�◼�=�h��&����ȩ���O1�����V���17��q�]��`ψ��A��߼�����qbK605!?��-�'���/���`�;_k|�6=)T�Uݚ��;چd,�h?$�R�W��$Ґ��Č�N5��|믫<	7";<����h��t:�2n��aZՀa>@���P�p�m����~�뗙�A�@G�j�|��2���ru���_s����&���1�����ɩ+c�D�E�KH�'���Xo�W�(3q��B6]�u0����ꕅ�%��=�O��^����.="\	I@Dg� @B��DE�v	�<��܀�%��Agov%�S8Z����l/veB�Ij�SK�M�$� [�Tc�}���c䊶m���\A���޺C
8c�G1G١:i��>���捿J��2�@5�ۇ#
ύ�9�2�##*-z\os��ȖY�ч�5�#o�굘g76��g�i�A�I���Ŋd��G����Ӂ��Vćh�����bI���Z!;6s2B�P#��;4�x<>�JF��������l��Ǜ��yLiՔq,;`�,/J�ۊ���a�� �g���܃`\����h�&�|�n����$�B��m\��#������s��S&�8`9g:�A�`:��=y	���A�c��y����?���d�O+
���}�?����0Z� �	�@��v��qNe��1 ��p����yW�Ht��
�t�!��ώ�D��ѱ�"��fn����H<�����KU4z�{D��w��j�I��Q���_�����
'�~�<�$-��<3a��P�bԡca�`��fx���\��b>}G��x�w���O3�L���������[7��s�3�0/�Z��фj(ó8��4���4�rzU��B˘-����n��_q������:��n�w+�x~�m��D&!�,��4�l$a��
�Ғ<�����♏�"ƅ"�W�!"&+�|=}1Ph���,������g*L��5���M�����=�,p�:1�iU����"U�Gєt���*?����y�s��=��ѝ�0�Y&��lt(�B�0� k%����H)'��3����(���\��9���أ��`{�+����eȋ�ڹf[��D~A�e2)Κ� #��������h� �t� #���^*f��B�*=_�4�t�R6�Ϛ=@���d�뭣4}��_���V`&��;&����^�:�׈`�I����[
���*�$����a����NJ�Y�d�g#~��A(�	���{�A?�k�8u-������Z����~c̹1|է+_
H�P2㊷ǲQ��'#�Q�'kw��,|×��4�@��0��x��(�#��A�3����A��̩�~�vz�7���*y,���H�i��ĹX��'f��.=܀�vD.��#�zA�0d��Ey��J��&M�-��"-��ѵ�m��717��ߩɈs�Z3�0䓞����7tƓ�d���Fͷ{���$��$h����}ǛM@����K��x(y={&�FP���C'1]������.t�nt���kɧfR��@|6��Jyvc/�4�<����~�AΟ��\W��o��U�Ƴ��ov�p=�)'�I��ߚ����Ȏ�Sά:���*��J��D�8�wN��Ԋ�������)�^\�J�6\�8�"�

���Nsj����� �ld(&��ǌ7����c�oXߋw�k�"�x��c�^�k�=;n�
��f������}taLO�E�[�D�zݎ��L���5j�8w���s*�;M����iR�ë�7K����xJ���1�7���~��$fˮ�%�����]�d��al!���� OM�&*�)I��<�h�{h ȑa���t��>"暺�o�$ѕ��Y������*�U�T�7�h�A���~�Uz_~�0�0�h21�h\t����*�1�[���,����!�=�۶���<���ib���C��z�8l��$n5كC��/n�B1�Z�YB �W����*�۳�������A��P4��Y�����0������4,d���Q;lZ�J|�C�"��l�8,��F���N 3����8��h����L[i	�0��ǔ]����`N̩�/�����TkE3�㜱��f���S���l�I���N��� �$�aL�x�U����b|Br��M;tT���_9�L�?�jm3xo�+�M�k������s�,�S'�\.-�z����65�����XJ�d9����z��x�ꐔS���{�XXx%]�\!Sv���P�k�
}@#�-.H,�q��	+S�If\8�-����gE��"���v�6Q��z�$[V0>Z;�G�T[%A�L��Z�^�9�:HPbeISf�/ӱ^/����딚ғ�R(h�3:8���N_}����䁗T=�n�ծO���J1#���C��,x��cq�>[z�NKݒ�h��LAX���s��`�E
�+R��G�\�����ˣ�,�'^��i1�FJ����E����̹��]G#��s���|\p���n��;�_�[wk1)�k�9�!�KLy�[h���#�z:�|
�t�5.���ߴ?F
'l~O��4����O����Ov2A��W��2
^<ܤ������[�;����9���-���=�(���Y��J�֭�����4z��A'7^�L���|���Q�+����F
�2%m}=Q��'��k��G��ܯ�գB:��z�k��k��q�e���cn��v}�*��m�L �e�c����xk���?�)����n���%$)ʕʢs��b�/E��A��R��@�7��!z� ����`L໣9t��<�l���r��9	�1�ΠӈX��jÙ�	�f��`���35|���|�*���LJ�.�xc���� f�����WQ���v/I��~�GFo�gŎ��^���ùj���p���u�7�.��L4�Ț~�"�!,�0���V$FDכVl��_��@>.�7��e�ꝇT�TV�T��9� ��O#yI9t��}#�L�8�Ȭ�ѾF���;0��\Tfh�l|B	OS�؞m�:t虴АR��i�֝XWI����̊�ӊx���WxGGB�v�\:mZ���C��Y炕%#��sA&���0�7,�Ue�汮�}���Ц�?�X6K��#�]���z$p p�l �X�����B���r��Kq#��dî�r+ȸ��D�O���H��W&�~�J��M�%�$�m�Z��'���x�m�]Uqsr��&��ms��W�XL�U�{��&)�d����c��=������V��%ೢ��K�/d��ۀe>�;o_���������'�`��0SIGE'p�&[YNW)ή��Ľ�ɚ�^i>r�T�6Q���/"|�q���B</�{��Ե�١c>8��]R�Xo>,�z�*�s�8🺻�3w���@���v�����N��k�'xqk��r$l�ߏ7〔�)�=;�7������u e�j����W�.���� 3�������;K���$��#A��@O�F�]��V�:h�v:ǔ��]p(s���]i���!�F�*3�c��x�.��N���8�{nR��ݓ����J���S��*l�������E<����5�ʜ�m���{i)�������ϐovE@���o��	�Qr9Bn�\`# $˲(��X�EU>�w�ʦ����t�\p���W�ܾ8�����w)��7�Cgg[�h��"$%���˂���\�� Ο�}vG�7[�9_�y�.�C��q��>��� �)�2� �\H�)l��C!�U�q�6�m_�>���������.�^ه������d7��2DB*u��:{�4G��^Ӵ]L��&8|�����D��$���� z_0:P,D�9g��d%���UlCL��}!�O��bq���&�I+ �g �U��Sj��aE%�<�X�"_��L���9j�a����t0o����}ͷq���~!	�]��PF%�;��Ԡv���#�'�ҥJ7D���`��g�!� ���Z�jD�c�`rU�*��e�F=���F=Rq��ɧڜ?�TQ�P�3"�m�p�)�x|�|@�3��8���f*�7�t�%�4N�~��ժ�bQ��NB7I�WT��*J�?ш��BZ���������quzr~DF&f�M�����#r��<��z�r��`F�)�+� g��]��y\3�u��GE?/�����o}+=�������G�������Wo+�Y��᎙=�ykh�w���8��R)G ���`G5qd�8������/�Z��92`M{y��&��.��0���jRDS�-Ρ<�b<+N�{ӊf�9�J�ؐ��~��Dq���\e���}0���� ���M���7��S�x����V�|�GK�����I���d#:F�Lf�`����;e��b��RI����s��@����r��cz��<�']�۲tV���c��`@Zg����Ek���8'θ��a��o˂@�R�f>�(q���3e�G^����3�F�/���.�}[ZȽ��P�筁������No�;���B4�j�B����'�0`�W'΄�x�<���$'�4N��8����nx�"��+�h�Ө����z����A��=�,��졺���qY�R�
wVZ��T<σީ;�H7G��������OW�j������f�Z�A��@P���B���e�{��5މ�'MT��[Smb�K���gт��������_A��Ͽ���;9�\�P9�0�d^�R��FH�*��	PU$,���mEg&��q&���������*���D��GtPȄ�d	tt��/�m�͎�r}:y}�~dh��l��)3��?*Ӧ��: c�Y��R-�@R㰪Wv���'�G�j�.�O�̦�V�Ff�0vM�2܍� ��^�R-�c�u~��K�{1�6�hf���~�9D!�)� �p��Sh���5rk[�����ww/'����_ͲOqD01�1�8v�[+�"[��,�"ћ��B��)�P�i�^�@D�5c,0�p%���՛�˾I����$5L�Cʏ(�	�Q��ў���Rr�H��^(����'�p��1y�EHP�ǋ�^����7��+�e���F���o^Jr�BL)���l�63$\��\�e5��V����|A�-�N�]�PhvF.>(--�^������n4����<��$ƛ�TrxBv�\�bxMn�7�c�&t#�1�?��[S�
<���_��=H��j���Gbqoe3�@���p���#),V(EU��2��v["(�&Ξ��~1�n��Px�S�?~��D����
��de�:���`��"�N�*~RWP�_E����䶤Ϸ���F�1��!�M�A�������^;�K�AR�e]���)r-!r�ߣ�5��4d��=���B~� ��"(����C<(%�h�e)*WK�����Φ�fx���<=�jV2�Mp[��0: 7�_(W�@�={�51у)Ӣ�Ӌ��ŕvݴ#`�������ט��p�rUvS�4�~a���C�
�'��C )d��F�?�;�9��ﺽ2���j�0�����g�� (6M%79�	L�3#���Jl�C;�b�&>���M���3�7ſ���o�|O�B�����x\n�;���.����(��%Y���u����.g�}F7�����%nֲgI!����q�������|��	4.a�V.Ŗ�� Xbeɍ��J�s�t E�YԞ�;�F�;$��F�R$���k0���f��+@v5�[gA�U��7�:AA=��a0'/lBA���2�$�jz�:��O�a3 ^��b>X%�37��~�!!&GS�:w���n���$3��$�J$/&1z��13���e��;�@�k�N�$4#G�-��W�e�DOm��t���������z.� ����ꠁw�	��o-�ajM�	|Q�f9a��j���Kb��A\��Ԩ�&�ť�a���R�P����K�tOA�}פ�w��6:�><(D��w?�L����E�-1�d��g�;�R�sJ�i5.�)6߆�p-epF��yL��Cś�$*2>=Qt������a�iQ�j6��T@���9�]I���a���Ȼ����v��}N���a�r�v�o�k���ʹ�I�8w�x���N��x[�tڹL��8Xh��\d�7*�K7��s���a��a�����=VH�,o��{G[�K���:�9�M`�����������D���0�d-5��ʖg�%�v���`M����%t�J:
����j�:~��c��%xp{7��ɻqh�9Y��<>ng�h5�ɠ�R�7=I��n+27�{��?60>��h��B<_wp9���#����7Ŧ�:`	�Gp�ͤ���"3"Fj3��=���\�g�{���oRΜ� �lj5!���k�]M�NF�uN���2Ѐ ۻ�/�Khjг���7vє��t��W4��������r~���V�	��e���ǔc�0��W���� �l�0=�pѕ+��N�.��ϜB����³��/�?�V�?~��F����'�^��/Ώ4���e\�m���/��C��YEҹr����8��I�"Y���d���i�^�H�E�5� .��,V��rx�D�Aw�6��J��\����򼞖:��T�LX�V�0]U�	�o0�-m�<�]С.��4������A���~_�s�y�I+8�5�͏�����ؠ�&s3�"d0%E����\%j\)�9#W�҉kb��-R9��?`^��rm��m����ԅ�ҍ&O����5��t�,t̀�o��X�R���j�N"x(��
s�'S�4$E�b������m�K���ђEj�q��A2��������e�FA�}.�<�i	��c�����_ұ�p9c��C�T�>K5����Ŵ�Y�d5��)$�8/��> ��*��Ū��Ǡ���k":�ߦ{ZR@QL����$��.���L�$��"�&1�w^�1}HF��޷+O�!�W��K��a�<�A��^����*���(:���.��v2�y9Z��J��>Y={[;Q��Z�/���Ʃn�� ,Ua���_Ju���b��j�<������_&��&e�Yo�5�{�⾮�������O�@"d�[�� �O��O��Q��z�U�TO�v*$��eם��nb*���8��G�|v�{���ly&��@��3r�bQ4���U��D��iu{3�ث=/�Ǯ���e��%�Ą��ڙ1RܻcG3���dD�-T*��rPC�Dv�� bi((����R ��m��T۔YK3@,�a �ڝ��� 򶻁�P�3����4Qx�כ}�� ���;�.Z5Ϣ�
k�垼�ቦΰ��V������ﾠ����q������P�F���`�=]��3�{�鴆��f$(�9�8�V{29KV:�ɇ��ѣ����dp���qI1<ű�zi� ���
����Sz���R�5���������T<k��)�dK���=-���=�.�9�~�;k/XA/��8��R��bs�.��L����Dh� ���dnf�����7�`j'�O����4\�I�N��������!��-;<"����y͝v��(gY������a�6d$d��"i����2LI%g���2e^��بK�J;Txd�h]?a��}?�Fr�-��s�̔+_���J��L<��|	푱qlpy>3$��;d�Dj)i3������{�^3���$�M���Id�݅J�E*���Cs�qC_$BQ�T�Ǉ�&�����Ψ�d��H\1�J�̓h	o�\K�[.��aԍ�{șfp]C"��ޯ���M�i�`0K[�3\_�HG$MS�n����ym�
\n�sA�XU����qa��,����;�NY���<kg���c�w�!,�L�!�t�bj��ձ���y=��������,�0����f���~7B�+����Y�K�D��6��EH�/1O�1�H�6e����nN9R�C�0��0ٿ���:`o:��|��3�N'�&4��D���ì�Q��uF�,I�4�v
����Z/����.�����n���2��6A':_����	�oQ��6��Ua#H����@��s�"�{������e�*��md�Y�V����ӌ��!T!!�����2�������=�3W�%�-;�m.;V�!����l���-�QQ*��]��hS�%�"Ѡ��R�ƣ�&���#��p�ਗ਼��̒+�YE;�TD[r�o����z���Ov~gD	�����*昳���7�ʮG*;'P���$ ?w�5g��B�A� LġS%�d�qK��9�=f��K���鼽(��AF�^t>���и��3����D^���kc/
IE,k?�-�+��Q	�!x[[ÿ�xM�� �F1�y|�h>�jK�en�u;pA@v>+{szM���߲Qc�B*�$�cR��"k(��U*��ƒ�6
a$�i���3n3c�S7���S�?�uf�m��2C�����N����0ȡk�h3k�1n�#���L���βg@U�:�2@ƴ�H�j�.N���T���r�\R���gm���k�B�)�J���3!�l�V����lJ����zu>�$����4��Ǖ0���%�L�S/� ��8"Ԗ�lC���tUʐИ<�x0�f�p�M���%=0m҃�'m$a09W!n����պ_l��+�s1�^Y@���/����z��]�򠠍,=���Z�����!n�-ǩ0P�+�]Bjo4;	�sD"���B�+��7e�>�:�����@�R�B^�����mDz~��[�W�?�ֵ�\��	������+x HJ���OK�2���5�җ*��c{�'۴�Z)�)���I?Ջ]�f��=�K	�,�xL�	.gZ�O��`�%y������,v�%�Q��"����=��֭���d��N�@�����?��Z8B�A��y��p�u�yr[ηV���h���U�/��U�s�F���]+�w��Bg��S|�lR�I}� ���j`������}8?�>��5_.��=�P|�
���ǭ^{2���H3��i�i�<V��`��3�o�+p��K��ѭ;|�����#�։��`8�F+�a�)���"S������m�	Osf;!�Eͽ���y:Pl����gY���#�N��a"�B���T7�e���Y�����d��j��<U�;3x�a�:*.:�����$Xd3y:�� 赗��v0/C��<�����{���'1 D�iƸ�Y^���m���J�3�kN��b9& �6���L������!_����x��w쵑������ ���C��Y�'�d0EJ�~8�#�ab3�;@xm�C��eKf4�2��Y��Ȱ�������ơ�(e�s"�xh���z;���_N�r�r�l�����A|��ܚb1B"]Dw�&J�U�R������d,g/Sd���ݤ�
)���M�BƟn�@[[mr�����#�P;5���H)�{�I	�h�1D�J��w�� ��\����i���-ܳ+GYG3k��_�XٳFF��^�@�;�!��(]����ױ�c�&�����M�C�x�7�=s��~����pI�/�1�>Eiz�/��.�dDC�|��H�|��s��],wm�{|�������5b��TՖ#�fҥ<�8Ӛ@���4A'�@�;�Q��:�BKt�7ku�
������m��:_�f p"wiy�a޹�Q�߱~
2���d{q��}:�sܩ�@�������GK,�qᖺ�R��+���&nQL��;�Bs���(2
A)�@n��́`MuZB-��S=B�X�W:y��~�����̒Xx���w]��-GT���'��"�LEL�I^nOކ�FE�b"����{�1��[�
D'�R��Y!�_�&��]O�9z�o���>�K��Z��
���Qm��PM���س��D D��)�$�X����[�JTk3�gA�?z|_�V�j?��k@U7�߫�^5c��2*ػ�]Ԟ���i2e#Nk,��jj �9�����X�J�ԾT�xi1�6[�LG �"C���7��8�::��?���W��wۚ��=&ڗ��B�l!��o�q
��c7�AK�TEX!�uz�I�k9��sKM����b 3�V\ѬIP5����&=q	,O�}4�~���پ�L��0���I�eq��!���
x\9Xy���)Vf�;̼��[�\ѵ�o=��|O9/g]P�l:�+���-�]��r�B�^�[>f�^\!`��	Nl49�#,L��G��XWL$Kb<����E�H ��_�t1��䄠?����ȩΩ?
Y��-��u>�?���K�i�	
=o���H��N Wf��I䲇�J����d��_�
��q���ۭ/;�w���1?7��>��j"�8�(,�a9�P���Z쥏�0Ȯ�n���BO�ױf��J����k{���pOEBt��	> � �k��b�5�����rز{U�� �v%4� ��?��ow� O{/u�t�.�Q|�E�F�U>�s������<�#�(-�����Pȱ���y]}>����<+ -���9�����B1�\6�&h�CÜ��״䕃��}�'B�1Y�Q7�Sm�3������������<��P�{G�{�^A�h�?s�q�Nd�c��Bg�Ba������+5�y�4��;��6.C�we-{�J�N�NW!��C��1�?�����!ֶ�;$��B�ˎ�ZN�BK.՚Z��o(o�(�{/^'�ej^&�����ߊ��+>Qv%���]N�[[���k�$�~��`�E�r��rx���W�D��F/F��� ��*ʁI&���fB��tfra��ʀ/*�HV�$�d�T56usu��-|`�x�B_@P?��^�zl2O�#��X���M�y�t����@�&<�*�wPѩ���I3y��j����/k�j l�oi)q�j�i*!�\B��t9��XH����UD(�lց�<XYh�Kn�� �� +C����	F4�l��\�c���mJ��Y�m8r���O	����s����i�><'�S��nbR�a��Nl���LZ1=F(f�J�p3�i+u�$2�uU������H,Y�Lcd�ݟ�)5����[�����]2�;݀W��g�2<xuZ��!�k�j�S���Rlß'�%X�נ�be��AP����H�I�d�d���}�+�9TX���;�(�tW��hzԒ�aE��"e��S�C$�����UH�U���̾���}õB�� �ۘu\�7�!X�l���w%�vA�Cd��ہС�L�,��N�/.��,�&�3F�gC?��W�U�٧�-����C�D£	*2e�D���dE3�m�����l��r�[�=�	=�
�$B��d����Vi�,)_�D�
�8D'/_:�ƶ"r����W�
9�R��<��oK����٪�h��)G"gV���:@=�����D�����@j"��^���-� t6�ϘS�9���th�̜���y�D�����i����8����:@I���WO���5��s�R�nC��f)`�y�PȨo_���(�}}���L��
�� ���'uιo�@Nvƴ�����;�
�\8�Aj�<����'����F���Lͣ����at����\ʷG�&���'x�S&9Pֲ�VZ�0/i�ɂ#|SbJO��M�P+���OV�ˣ
���&񑛭
�ې�o5\ֺ�&2B��|!T����V��W9H�&�ʊ�	5��xo1�W���_υx��j=Mj�[c��b ����񾲭�@t�J�:���=��s�s}/��n�K,b�ˣE�3oY5�H��*5O͓&�GP�����`VFw�m��x�^�l��[[᯷�g��!�b�榗�����~�i�Dg�0��
��vF�ۉE3	1��r��Wt��A�[��lm��9�:����<m爐�%2.,~|(����C!�_�����K_s�}�g�~�{K[N��Wfq�Wu��,�B�8"�7��)C.��1!�u�V�nhՎ	e1� ��_��JK�(�aU��-
�\�n��IgO���K����8��!O�>x���v�Tt�*2�puHy`�[R����Q��Lí8� /\�nk�L{;���th��j�(*GQ]n()�9!�X���Op�P������VSk+}�,�^�]��c�w�M��|ӻ��Uzt,�\�h�X��Rv�����D�X��վ�s��ِ���y�u��.�@<%�'C�[t.���ۿB�}1���'��R_�J�G���g3{a��|7sYV
?�=if0����+Q�W�r����>�9�_}-*���#���� M�LUS�z]aKMZ��'�s[�.%��P.�F�.u�'��� �?��iu���0�K���86!(��%�������@���aq��5����_��9����� ��q5���\��Tk(��a�]��R�a�x7/w!KL�סG>D�|�z�F3�����Iv����5�<��˛�d_����Xz����$#�`',��v�a���������Cf4;E3�u���_�s�^^�J��AW&ceA�o	��@Vn���N�zĥ)���p��5cxݼ<�N���a7�b"n�ȟ�[���T��d3��V3��=i��2�J$6[��x(�y1����b<ͼ��`/[�����	����F�ѣ�C�lX)�u*��3{�����OJ4��ܲ�gN��3� OF��A�:������+g�W���Jʉ�"b���Y3�"�i^�z���B5�T�2�Kg��r��%�ѿ�n�c��:B�lE&u������^?�k���u�ޱITE�{j��\���sn.�q.�����Z]�1���q��
��Z;�FZ�����pN��gB������1$��$"��7�*,,��LL�)Q�&D@�O:�4������I���*��N������/�N�ڴ!E�U� z��.o7��n���{���6�'����<v�_K��"Pa�t�sw�#!�'B"��o���=����Qş\�B7\� #!%��ͺ�yZ�}�TCJ���*��������Ś�w���n��0�ƌ"���hZ`�g�n]�1Zً� 2@Ϳ!Lᮻ����i]�x��"�b	�ѐ� �����P���J�fs�^Es�b:���!L��H�ݹ��U���SR�*.t��{D&�,���w���ۄ��}���3b5���Ǭ^���,���#�����x�7��g���-���j���@s{L�V��%<��8�K��E��­�#t��S����g�s����Ivr���@����$ � b,/V�msN�]>!��rn���ա�Ӱ�<�˫ &xx8f�jl8a-v�vIX������=bi[tu8VM�s0o�804��3L�=��m0�-��*��3�p�x�,�}�5��t
�BF�:&�J��[��J��^�*����;t���K��}h")n�Z�L����8����b�z���I�58Ї�濈);ᎶV���Ҍ�x3c����@�]�h�C@�^U1�ҙ���ah|
Ū���:���S�Dxm�>|����?2&�"g��j_���=@���p�B�g.p�P�M���UG���b��N)b�s�t�
���:!��(&�6�~�\�ABa_&瑞K�P�F�Q�T���1x���b�����D?���Zx�����1�A���l�\5p�kR$s��L�LF�����%��`�ν��N
y���|�|\��ؿk~���br|XH��t1��`$�Z�����w�u�[�
�>�ߋm�����zT��tXר�_@�G�:t�D�2J3 ����YE"ڶb��;��<gu��i�g���{�n�ں�]�n�=�{\��V��f8;�lW*N	 !�EUQ�&GJ� �얢q��(��slk�
��'�w�H������ѸT����
Gc������p$R
�eEA^U���ᢠy�����IV{�L]��C��h4�S�`/_�f�Xoj��C�7��ť�͈7���n����i	l (�{Y�مmm2�f&�D�A�g�:V^�{v����T�M����C)�s�Zq�'?�ŋ�0�*໷���GE�B�4ڢz
"����p�2����@���B{w�Ə~rz�䆥����}L�Ag{�����C�P�!��� 9����0��Ɛ��D&9)�f�u2����Ѩ����-�h#��Z�����lݵ;�`�!��%+�c��p��5��Դ���^xv�;��G��=�U�ף���<�/|�s�Jg=��Ճ���?b�	b8�#�����	֎+Ɉ�[ǧ5�m٥�ؽ
�.���;� ���.�d��|&]󐚚�SLCsK�TGx-�0���L�����Z��K�@Sm��9�l߹�CP�l�B0ކ�M'�&6�jyOG8ބh��'UI�b|m�\^�?��HS�:�őpzzRFŚL&���l�[�ל�t��sYذk��tJ�� �n���bp��cpם?�H_,Cp>�3d���������?K�Nv}"��e��x�\�Z��p��ٌ�s�vpzc�L�d����TO?�
�3ƚc��'���X⟿����d6"G��sK�Hb�eNb�#Iy�[�1v��	���ŊE�qԑ�p��eHD#`������s�M.�X�JE�k���9�����siijB0���Z)�S5?���06��+��D��1?*s
e�<�(���,j���Ɂ�W��td3M�֑��{�����{.��,]Ȇ��y�gKY��(z�'�e�aǇs�[q�'>��}{�y�s���_`U�u����Aȯ�<u?H�f�J[��g�ĳ��=���{}���+�z�	n��sOK[݊Jz$ccl�4��/,^2�G._��9�;�6�y_�_�'{��q���V&&o*��� �Y0o�bW�1J�뤗x�Z�w-� ���c1�ڻhm���'Ȯ=�T� �X��#���b������ő�/�Y
A��)�&,��lـiyJUɻ�K��bUEJӴ]3�����d&�P��JWU7����S(UdU0��ab6��d
��Ķ��Ѐ��f�54 ��HOO®�D�26=)�HǼy蚻 �d	�>�	�v�ʛ7K1�FH�0����,^؉�T�����qh E��F��=���W3��۸W�݈h���8~��o�ē� ��B�t�M��{ߍ�]r":w�����`b �t!���v��A}����9�e'M�KuxP�A��D���V���L=��ux�����&B�1w�B�8�H,[~$ҳE��JQ�EG4���|
��D#-��E0d��K�������Q|��M�]��ނ���R�"�'`�d5�'�1)>�J��IH��	�r��Q4#QX����&��tK%)��R��,,ݓC������m	440Ζ:�u��:͊��0�&T��kN��DWF2%�KI�$.�YV�8|E�1����b�d����1"ҥ{�G����r-,���R�QA53�F5�37�D<����1��z�`�:ο�\t�C���Ǎ7�(q���t4�#(�2r%�`%S7z1��}��H�.�-�H5�}�E��׈������ַo���_첳&�G��%L�*E��T�f�2�jmlD.�0<���Xu�2���@(`!���`o���19=%�w�P�#��~��5�g�	��Ʒ���s碥��'ϩfRYI�-}o����:����B�"�Zl��0'42����L<�	�˘[�]��֯GCЂ�9���`�����#�$�������(Uv�t���ڄ�|��:t�?�0f&'�Z%ӟ�)�q>�3U�?o�s��'����s��$��X�q�r���	��q���}��/����H����y�x.�`����ɤ�k����B���<��;^0蹮뙦�ض�+���4%Q�>n������R0�����C��,����r٭V�^�\�J���6��p�u�.�a;�y���Y��z}��?��_�=�3���^���n��k72y�B.�4�;b�H&�$�P��PZE�g�:�Pzc�X��ؖ�E8��2�<�G����yA���#���QP�!���8���V� �.R,�Le�E�P��k��+JF�6�)�~M�vUu����s`NSM+h���.yPg�U�h\a��X�7�У�5�kh�E��L#���`a�I����)��]#x�׏`۫��
a��h�����]���19[�w~xv�CA!�A���s�x�g�ӎ��8�{q������aL�z������p��ލ��!^��������u`r|#�����Ĩ �ej�[J\c��E�5��Ѧv,9�hNe�?��k�#�y�E�BQQil��EK�hl�]�	Y�@SX���f������'�A(G��<hkV/���%D��x�7����,Զ#�F�����$|nd9Kg*^�����E�/Iq:�r�%��]��UG��r��6�"���,���[ _� ���FIb$l"H_]�م 	J�=�#G	���Km���ds�$�����������U��f��˵4qdaư�������:p8�$�Й�?�ߑ�=��Dfi�L?����Л���'�c�p/�F��\r	N;�t455���ø��w�� _:�#�<�c<��Ν��|��RIư��v�D6_��������O?�}��rO8؃��t�/�cgN_����&�y5�:?[����U&�����S6�!E4��������ߏ��)�R�E�?6�	�r&�R��n����Ӧ��{sk���r5���%L�\�,d�щI���+��ۋ"���DUg<�*�e���_63�y/)��Q�<�]���ZcQs�G�Ν���:G�Z�"���3x�� ����:�Js����/��{�~�:�So��D@ 'q��[?�*�����L��3g���;��=�1�)�0>6,	w��,Je2]h=@)�U��u����`U�,��p'�էzڬ�i����zj
򊢑�T�H���UU��N�'}���ӓ� oq��<�Vu%��L+��3)�
*�Br���dш�SQ\�S���+��+@՝YQ�"��k�4����t��tWU5�UUWqU�S=#`8:���y�g{��UOS]�0T�qGQ5��tUU�S�?2�UOU]SS��C��V����N�=�寿�Ou���~cϖ-�#�� f�mU0H�����f<$i_rA�&B�8��L��t�(щFE�]R4�*r�����czjV�@�1�,C��܈<P��jZ��MS����Lð�U��+���̀NtvU��c{Mw�V��\�6BΑ�ˌ��>:`E�2��@g�7s�Ɛ�|�5��TG1!�ף�b�����7H*S���0|�^޺���¦�c�d5���|��X���6�s���g9����uKu1�1�+.9g�\�`^yy��o���d�fɈ���y2>pٻ��E�#J�M����,�]`rl��C�*�F29N�	�3��C��u3
6�:��:�x�j�O�1�*bہ~�������xV�=�B�398�����Y<O>�0~����XaM�Xҁ���WikƎ�,���O ��x��-L�\8eߕK�e� ���<�M��:�G�V>IG������IJ�a�Cr��oW(��������FBF~L�BR�����F��BO��!��!>��"�T�^�+�aྖ O;X���9�"�UN8�61'nl��z}��F�N�%}��c-��(>˽�D��@oin@�;,�2��e�]"z"�(���Ȉ��$X��6��4����6'KQ���JF�@0$������4%	��s����8��o��/>	��L�T#�͏�+YNUw�\ilQl�<�x��Ւ��A<� �={�K�#v�U0�.����rGNFX�����>��пf��W�+��}���X�h��^4_:�?�?<�<���B�[͐��k�9�v��E��Y�ܫ�C�����z����`�����W �`�k����-ؼ����F��y�����؀�_� �����)�Й��뇯����|~>bU3��s��³���9� ��׿���uu�)j<49���A�L�a�ף/�S��AYq�æ� o���Q��7���'uҝH�j�"�h���|ԭy��!�����ǩ=��&�G��7�g����{*���������/݀JF5�<rU�J�'�h����O��&i�c��~��(���;+�h��*�gW�
4����`$�s~K���c������������Ɂ�U	(����(�aswkS���T�&�w!!��K�*���Xf�g����v\�m[�z��#rAҕ�*?T�/	��hd�u�x"}�Z}���X8{^ūTX�U�R�ī��Z�R�غ�T���f�F����u�eG�˕9%�m/�'j�Aa�W�iJD�"DJ�x�S��q.�G�Ñ8��FT*L�
�Nt4��x�l��g7m��/�(���W���?��X��c�6�}���Y䊁]3�Ґ��9�ኋϏݷ    IDAT�y'�؟vp[_�&���Ff�xg�v>��K���EA��o<��}1d��tzr��)LO�H��ڲ[����E]c;�J�cŮ��h�jN��g`/���D(��F4�[���bp����YS3h
��>�֐���0���S�]�S�҅����B�	l��[w=�Ē�1�b&��fK�/����H ������jv]�;9����7��E��rEAnfF��
��-D��C�,*d��ޓ9��X@�$e���Z3M�vu��O�\�l*�b&dsŢH4�H�^:���s�CS��
�~�N[�E^�����DI6{�Cg�O}�.D2�c�7 ���R|�cnRv����g?����\��EcWF@�Fb�z�O�
�Z���H%��q������IWb�S�֢>]I)�c�C"Y$����_ݎ������dJ�I?G�ײ3������ɉ�RaIcPE@�|��}�2Sȧe����`|�/Dx�p�`0��X9G�5��:��YB��' J��q*	G�9��&�r�j,]�LCW�B��Ŧ-��34,[�ܩ�'���h�;i��v�����,�7��U&�XX�Չ36��ǯG�0�i��x~Ӌ��NF0�͋�4�t�J�8����������:�p���>��d�^'�����s�N0'g��v6E+W�ĥ�^*^��{C~��rF��K����B�iX���{�3A�N0
I�����|Y���~�|��W����e��/Af�L�����:��gD��R���WD_���'���_��u��ڏ�F�<�yD�1�Wy�ձp�}��X�,e����tq	����"۶�X,�y��E�-^�����֥�����w�穓��t�-[��
�:HXS9��o�@$�ZU���Z�U��aY�;G�⻄|6��|Aؽ�&��,MMxCq�70()���V�o�q�Y��=k�m�5l�vtL���ׁ���Xv����;�g�����nr6�D˰$x��� �J�&����{^uh���� O��w���H4�Y&Y.!U,A	�p�p?y�w��M��Gએ~�V/��T	���`w�0ʺ)��\t�KG\wqŻ����>^a�����;�C2�F ��)d8������ۅ�H�8��tۢ8 c����^w��F*9��� :=�i_K9�}�0���t���Y��)�p{������Ζ`�0k�X��,\�#�(���h�RJ�+a"��QI����=�b� �������g�ښ��'��}	V�j����8(�b�N�w	c2a# ���?��x3�����(�{����ζ
�P�W�K��	�^}�����Kg��#n���h��Q�¥�`��~�d��k�J��Դ�3X�67#���P,��I���-�U���bɟ�h���:F��@�M?��G���������$?�E�I��u�	�q�������~���>��r=�]�V����ͦX���yH���]�m�()����9�)��AV�
1��m�b��y�6��׏�N��D<e���Z��R��aP4�4�X<_���vw��<�Jb��ػ�51c�{�b����y�F=��'���_�{�����eI_���{Ir��*,�倇�ŋ�bŲ�X�d)�+��9��^܂��u2���L*��7�%����rO���̐�2�uG�ĥ睋���I�Mrf۷oG�P��,[��Q�6���=�p�D3��K7|�vn�c��J����Ȑ�k�ȝ�'���Q&)5�F��q����(1��:��������&73)J�ёdӳr������|��k��Wp�o�_���e�.�Rb����g᜘�FZlykV����Vi��������7�豈��Ss ���_�_/4�Tc���oj?�͏�{W|����od��r��UP���˼>��.^��e��<�)����{�YY�������i�3C�*("
*�"(*��5n�M_Kb�M�����w�&�d�YMb�����FT�X����vz{����}��M��>���]�9��8�9�y��������W����+t����l�t����-`Y��UU��`M�@��ػ��3c*���̃������)zl�+�4���Etjk[��F��Əo��7m����}��q��eqFl���7��W^��{��9�cb�D�Q���[(���Pա�Zf��_nj�|Z�nt=N?�C1����*j�!�9X�0�������PF�q��1�ꗾ�Y'OE{W��������!��b�P@��B��r�R\y���iӛ�ͯn������ޖ�s6�ⲋ1��NA�C:	۠�4*)t���z`/�z:��ٮ�;5��U�׍��z0,
���r�+�i\�M��}Gz���Պ��z���0P�b��騨�L���p�rC]�PGmȅ�_��O<��T�A9�SO9����SY��w��'�D�SqhЍ����c�jt̍���Nb�Tc�r̉�W���oC{���[|�\�  �\^���ɓ�����Eo&)�b�M����S�&ϓ�
b�̙��m�]B�@w��� �̚�@$�he�f���8��g>*ٱŬV$HS�K�K�
ȘdJ��˫�N_�B�>�FX���l�3�{���G�kK�:�P�w�f�<�9{d�<��M�
�|=G����)�4ǈYgS� ����Ҳ<����7�����s�7��B'�+��B*��SdJ�B���UQ��tf7�LJT�];wHَt&��ЩY��+Lb(�-��|UQ
sa>�4ދ<t��9�[���x-�L���� !U
��w�uk��j��*#��@i���t`Y�d�!��柆���]܊E	�Db���hg�-ǭ���+��a̟�Y��m���y�|�U<���2y"��nz�L%�>����0�-��9��^��@8���[�I�Ƞ��P6����8�v��H�)�e@����{��@#�C�
�\�0�x<��P��	�,�>��@o���]B�ʜ��s;��Dͩޝ �jY�2'�%�����Ȁ�������.�s//�S���k�SL���/��/��,�C�'L���N���ƫ�!�c(��z,�*� �r�tiGf�9t�xX2C�[�n�{z�^��yfS�1s*Q�+OiQ�f<�(e�������R]�xL����[�MZ��S�}c�ֳ8;=�����3O��Ic\�(L7���������C)K��!��J$Ԟ������<�k�_1�q=�э�{
m�ە���/	�̙���~��c��V��d�RF�,3�|w�,]��\|>�B@k[V�w/^��"�u�р������a\C�@q&%%�n��VZ[�!U�Ii��N��
���<U�L;�7��!���\ȖJh߂q�bOG���������NI�
W">��x5�A�X���u� �l|�q�:���^��V���Ӹ�s���x��ź�r�R(�{ �B֠�iZ" �@�9��x���4�_Ӫ��g�t����������lsZł�Ҩ؅Tц�|�L��C[{��u`h��-�%��#�I�\ġ�#���1���9��M���#T�@4^�L.�=��L�lcv-�|��#�Ts�>l��}�l��:UH�����G�����zq��y��]����6�@>�@0��
i�������L�O��m�usF�k[��z��϶4K�8��� �P�����Ѱ�l>7�9��{�����\���p������M�%�U���7"90�Q ����k���ť����L�h�P�2o�sH0��Э�����9�"9�Ԭy��g`�)��SZ��cضk��G�1�Ϊ�C?��IT���:���O��c��Z�D�[;
�lZ�5���5��r��N��u�~h;,-���n����ǿ��W^�㏮�!ۀ�$IP��~M`���TL� ?�N���̙#A&F|��x^0������VtiC&=$?Q�(o�Nmn�!u��ۦo\1��>�;�x�m/���˅`��
(�)N�\��x��<e�)w��ѶeY��zʔ�s��n��/��'t����d�v{K��E��-��ssR�v��.7���[yDx��kܝ?)�V*�	d4��3y���r��bҘj���u�[}��.��:I#��y��a-[�0��v�#��M���<���;�?Э
�P���*�lǚ���ά&8����ȪH��.�ev��+�缍�������`y��L�2��0���\ϡ`0����ڧ�U%n͛��Gn��ֱ?�N=N7��O��:��3����AM���DA7g[�B�ص{�2Ա��E6�#lf�e7�n?��wb�O��g@-ARe����;�x�8؉�x��/x�����~(��K�1m|#��5��do��
��?n4�R�j�\|�r�5�T4�m�6�E��E�������I--�8r�v�@6=�ޞtvAe"��.}�CD�S�6_@�"f�:��G�WV�a�d�f�x�@;^��>�ڱyO�p����?K7=��L8m����"��|���Iu1x=�u���1k6��~��ܵ���9���hΒ̚����J�#���d@7Y�َ���4 :F�ѲG�*t���/D���͉Ʀ�4�����I�V0[��� ���5o�X�[9�d�� "�L��s�����F�q��{4*��g����&y�2���S��0
�70�\j�{�� �5�(����x�U�"R�;��u R�����G�Ⱥ�ع�=�.�m���7�R������L���;l�"8��wn4���y!(��x�P��ѐ�芛Â��2
�5�<�o�r�%TD#��L�����a˾={̇��g��0�F�Jɡ�W^L��Ӵ�
�J�l�3���y��=�ɌI�B�F~|?��7u*�_~!j��0��bǮ�X���8�э�/����U�۞�&A�S�6H�tc�qS1{�T�زEI�ܹs��������� �B�9Lׄ����x��������!.3<���uŘ�r͘4�}r�A�Q8<<+g�v�<[ܙq-ٺ�9��cp��tҦ����P��D���P�Ȥ������'�_c�T��x���+�b��"���/�w�}>��[pәKKT,��e��������A��0����t���<4-
=�r�].���w��`._�K�>�_���|���)�U
J"7�Y�����^����r���f_�A���\|%𿋡b�q^�q3?��O����\.�K�+���b�#�HTl��f͚��qJ>j&�gYV�\.|�Y��F$����kk�%D�J��-�Ƌyeڬ�C�e�k����|����j�	s3��h�1�ݮ�H4������'��izw���<���m\� �L������'��C����)�0.E���Ԧz̜<�����ěooݨ���PX�>Z�(@�A��o��Ͼ��������k��y�N����r��vV0����Jp���x���[_�"fO+������~s�o�& �z���q��2�����<��ֻ2Q�SO=ɡ~l~�U�����S�"rzy33l�fWEaO�4�
����E��	h�@O� 5��;�!oy0jtb�
4�L����~��W�Rcjxp�x��W�Y���4�d|�_A���2��mk��ύ�λ])��?��PF��D�+�k j+1�o�Х,g]8�{Q�7(i��ۼk	V/�B�}�J`<?d�B4w1/��2��6���O�qߡ6�IAu��gFkf�(fD�Q��OT|�t
��_�ĥQ��U�x?���]T���
�l ]2�ଲD��n/�
�9T��u�'�w�,��D<���<�w����,��h<>�4%�"�V�"�-QJ�r-u��Ix3�%����<��R��Ov��CO�#�8���n7�� u�C�Xm"�p���[��Q�����G{k��9�lYMF(r�5�n��6�c�s[�@�D���}�a�5���z���S7�������}�bL�z�
�'3xr�F<��u����G�� ���[��1��Eb�R�Sƍ�_\z1fLl��n�FUV��.C Fw� SY�j=�G7<�}��3]!����oa�����uH�R��Tģ��3�`"��ɴ��ڡ��p�������u����r��M�N �2&@�
��d���$@x*�~�+;s���,\x��>{�9������s��M��匿���[�Vy6O����wo�_>����k��	�P�`Е��F"n&'��~���u�G�$ŗ��J+�͖B�ѣGg�\|�#�sв��&˲j��.���A�Pqd[D-<��ɜ�Ʉ��'nl1���l�'�/��+
�xX�:����Ʉ�������r���w<����GN���6u&F��ǺG��m����0�*�yӦ�)@yD��=G0��a�G!�.c�	���^��xCQܿ���}r3�Buu%���pq��?��Wز{/� ����b%°
J.9�\�b9*�^�^��<n��ϥ:F���3�c��H'��"o�7��>�V-X�s�lD��޵]b=l����e��%d�-l�	
#ҹ�F��͓��'���C�xo�~� :?��q3N�ĉ�Ma7 QW�%4#]]�_��F<��E"D+�������H� ����~y��cp�+П�)���:����F�����*�쿢t��SD:"�m�m��f�D���AG����5y �!L��|zy��`
��3�I
t_k��nݖ�|0���-	.`!�hs�y�A�׎nh���42ɔ�c�ٮ5q�T蚡���Nl ��Lx)ܤ�ƌ��V��J}��AxS����yb/����xs��ꜱk���ɑ�11 S����`G�ي�d:�$�&3;�w��1�F���b�s9Gv��,�A
CR\X%T�"�:a<.Xv"~����oذA{��'��<Ї�
^{ɘ� f�������M�vb�sv
%�R^Ke�}��������ƍk�i���q3�Wҽm�.�{�)iػ�Q$�U$8�Cm����X��� S碥�`Œ%x��xd�,Y��\~�|�m��uZ���[p��G��k���fPʥ1q�X|����;����Y���
�2����@RI��1akB|��a۽j<2t6�Q�xJv�Ώ�M`����SɻE����=���Bn�I�n�Բ%?���{�������q�@	Xb��,���q��j��������S��bF�Kkn�
�lV\.�sy� ��(kCC�����Om5�H4q1nL�x�g55���r�����0��v�����G1��Q�؀G���@q<pbn7f��G}ȏH9�@.)�MS����HW��f4���k���3�U��z�}+ї��[����Ѹd�r\|�
��~�7bӖmH�3�� �
"��yz1c�x|�3��)3&Hʵ�Hn��/����;������s��@&c�p�%�v�?���jk�P*%����f3�K��c�|^�)�o��l�K%*��<IV�Gzq��[-g��&MB��	�=�& ��"Q��&!�� ���;��3/>��׋E�/�g��ETWT��}mx��Mx`���LĴ�K��W��7��'*eU�E���0k)�� 7f�Fm�!��rh�fo��X}H,øjLAA��>;a��lZf6� �ǌy����#1^x\t�c`�d&��Y�#.x�DF��F�F	.��(�P(��������d�C��M��H���d�J��4p �|�,8U��ۈw����x������#�1����)���`N���{�d�ܝ�.@�g4����sg��i˳������E�2Dl{������؆:�cA�uaժUɲ��t�S��:I�G<�&Y�)ˈ�62�k�^*i�Y��bQ8����A�(�H\�������k��󓝓Ó_��Ͽ"H�JHSl(N��J$b�+�!�|�>�Ic���%�%1    IDAT��#���/�9�,�=�އ?l|��:	���'6��'�@>���K˘1���k���7��c� K�|����
���C_:]�Bh�V�H��T�V��1lq�eI�5V���);�2����Y�E�#w�T�1m���/Z���d�c����O9�G@����(� �4�p��a�=;�k�}����U�X��4$y�񊫚��N��U�9'�<l�3��T��r :��&���Q�o�\��c����u��k֬���y
|!L?�4�o�����杬.)�R��>DC<�ۅ����	I$vtvbTC=&�LB���x=�?Ё'�ۈ���gL6�2�嗬��_���>�����7�نQ���-7�n�
4	{]hU�e�-�K�C,�`d��w��]w݁�^}�Ǐǉ�/�n�G�ML��lA����#�)scc:4�gfl�>��`
٬9)PJ/�lx�D�{i��/��[�}����_>ge,¨��鐩�U�cy�����Hsh�>����0q�U�/��6n�gv�7�N_��7������E��wupSpeD@W���J��F::+\��T�}бu-/���8w�h����d��.[����f�a��9�|>l�@6o�*H�߶�ͻ�RcP��@0���f8^��<H{{��3��Z�&�1CޔSj�����&F)�(w:ą���Ё\����8�������ؾ�]��%���/�"�I}T37խ�d0�;���9��T۴!v@�?�IwP���i��@^C��]e���vs��C��Bèj|�k_��`$��֭[�~�z�~�'9�e`w��K�2GQ+��X��Hٞ�ˡ|X �t�5Y����"����d2=̷�C�rV�S&MV�y�$X� �پ���d�n�%�8.	`�� �R �&�W��sh���ݿ�z�t`���p��xr����[8i�\|��_�c�ã�=�r� �q���/{�o�3O=���>������p@g��������8A�i�;47'2��Y'���E
�d%�C��(�x�^���L�Lmn�cɢy��+�9�s���~p>���"Ά[}�
q���&5e�N0�x��K3��N�����h,�D�b�Zԑ���AI>�Y����E�R�"�jjb�p�"��r�Wo�2��5k���q�	'��	-�r�jikSa�T�"��2�ڰ�B�!/�bQ��ǐ$"��q���0vK��W6��w��W�&��XB��E����^�O_~����O���V9wѽ������-������0�:��.Z��.T;��?���yS���&rD��r�Q"��%��lZ�C� �M�6Ѱ�JZ_�(^TH�"��5�a��4��~��H��/R3(2�G�uOjL0ĠQ�!��������Ԣi3���y�c�S���ݵwܽ�x��hx�cƂ��W&=/��0NtJ�\��(��jrC�]�$Vbkҗ)3*MF��2m[K ��n4�ϔ�#&E���Jr�#(.�ϖ{	��q�isP�y�0FQ"j�S��'p�97�D�	Z3�'R�ҮE�K�Q���A�3Yd�E䨾H�2����$|���n���B����>�:v:��=Չ����m[��T�
�`Q���@I�F\1����p�.Y�9�N@?:�0�XӺ7]��S�s��D���̐�sg��� ���������cL�3'�;-c2���u4����'�%�.A��y���Ιh�#�yGV�1'$�R����;�4̟w�\����;�ġ�^�]>$y�Qh+���-�3iDxn��K.8��x"�|�E�|�=ģ��{��W�q�yK1a�4�~�J���K���$��n���ϣ��<����3��h�γ��8�������J�IlF��#G#+vg$���l+Y��!��~d9ZF᳅y.�"�Ǵ	��,]��;7\z�1���r��o|���=�5,k��R�+��� De��ug)��5��Ψ��J"C���HD��5��Ͷ�tǍ���1�yX{|�e��áu�"�k]��!dď���2�֕�W�=�uA'͚����X��!�>����u���R7
��P�
,��`K"a�J���7�M۶aO[;�$����� .[����Rt��'?�w���(�������h+�B,��U@fh sO>_��_aڔ�6U�8ҍg�z�vlGWg��F#<� m��GU�r9*b�Ԏg;qp0)P/(g��T�bW�����k��uM����`�������
�-�ߍh�U��d	�\!�'͝�N>	����"�:�����G�@�G)6��)�2o	�\���!�f������ˀ��L��
����Ht%#�SH?\��	f-:+�}�	�4 ;v$�Wv�V�c[*(*ZI���1�0�d����űX�Jl{��.��C�>?Y��r
�4?a�@�q�]nDb�H��[1���h}t�7j��m��"�DDv�v@���b�}+b�>t
"=������ۆ��	�i7v;լ�QP�/*�P܈��������3��S�a�y!��s´�MK�@8��G)VS�`lM%.\zF�T��"����b��U ,@ӿ��93�olX�x�H���5Q���eF
L��ȪөH�t'`��Gt�[�ǖW���!NN��#�PĘ1�b����(��x�g���1D�"��X)^QID�m�+�s�<�8,[�cG��L��ؑ+�TK6�˛��}>$����'�����W�p�܆��q䈸��f�̀.�Y�&�a���m�Ff|�5r����D�禺�O,&,yZ S��	T(�`4&�'A��S�5�Z6�7n���O�G�I�a_@w[7hVy��,��~�%��;�<�\V&��@Z���9q�M��BI�v�����M����R�4_ἆԕxt}$Vqm8n=�u[���i�ܻr������j�r�\L7>�Fm���кe��Vu>9�X���ۍ�X�dJ���(����H�\,!)��#q����������\���/���#�ɏ�m;�����*y#=XB��;��L�B�Ι����4&��� �EOgrh�� �=�����i�h"��HG�t.k�_��{�v�@GW�Z��:&�;���*���
��\�qM:P��'@v,�D��>{��0fL#r��$3���� �?B>���r�[��A�����@���"6�d����@-:Љr�C��;�^��c @#�'��Q��g�h�kt�*.�9;�y;�c�ߍ�������ce�Z$##������i��u���&"�ّB�04y��$��W^J�4���:�ݽ�F��4^Q%×!�w�hj��Ra�2ү�Uq�a���R�ba��/�!��`�mV?.Z�P�O?�4���*�^c��@]b�$r{,a�88�o�6�P�VS(�F���ٶ�.#5�$�=���ۭ^�ws��g�0nTV,;�rR�aӦW��'�ʛ�?�ωng �n:�g�[�<������I�@R&�����s{�H6�[�m��|W{�����?u��8�a�X����1K0*760a6�"U��nW��ô�͘;�D�kl��2i�e���=�x��W�����%�A��4�T�o�~-B76<�8�C�8��*�z���O���w��Z�l��:�`��p*x~V7�>s�{��%-�bQ)u
g�Aݱ�e��8��a�ئU�,:��_�₶c9�?y�W���~�r�~��������!�#�\EJ!��QE~�JR1^م��Bf"�
�Ɖ����8˔t��*?�HT]
����ͭ��z��U:��G+��B������J���Pϖ�R���_f��C��B���?j^Z(�c��ayi�b�=%���C������UW�ܳ��H?n��/��[�d�`y�P�����B��LZ��46b�f,Zx&f�h���`�pڂ|F���S�L6�h�����uH����W����oDGO?2���	?���x˘F|�keg��>?��o��>c��Ϧ%����P�ǥ�m��m�č_�f=^|�yͩ��0�.*F#?j*�.8��*d-$��`��:�)�� K�W�L�Σ�ҏ`�*����0��l�ٹ�GU�4;/4� �~�����:YA���
���g�$V( Q3
Mcǈ��74����L�(@:�NP��
�����u����ƶw�#�4z�x�\��9I�2I藈}c+����.r apD.�J!W
aw�@+�=�p��EH��x衇��[o{aS�����ǘ�H��6����i,#���P�Eɉ�(h�@I�3oKb�:��1�T�D�D�a1��� 0�*#򢹩+�,FuE�j*p�-�������7=�^{.`�ڑg��� ��T'��xe����hw'�i��7�AS�XIpMXx�(ߙ�(L��j˓����?a±8��s��~�G:A��`6w8��[N2���|�P5˱1/��-F �.C�<�Q�\,
Ll�Ƿ���엟�i���[(ds��7c����&W�� 8�|t�r��xu>�w�IikR��e�L�(�LgO�o�c0O�Bz.H|{���5lM,�qu�k/9��뮻r�1uN��L���؏'��X�u�p�����\w����@�dR)Q�B1Ӯ��Z�DU3{��ll�FR�*����D㱧����{�rWoz{��+Z���?=����ŋ�%��o��"`���P�T[�\jBNP���sI��$�he�(C�Ŕd���/~N�����q�/~����G��`�O	X%6��鐳��܍ ��&��'b�ɳ�2�N�d.=�Y6�j)4��N�]��%3wRq�3%W�n`�~��X��'�F oh�������W^)	�(�ר('�%�Ea'I��mZ�l�%i{J.7���,w��a���B����{�� �SN��9��"ח�tAܒ_/	WV�,V�)lb�;�?�!�`=l�IFXw�#v48/�4e2F�T���{v�Q5Lq�g�,�(E�т**I����h:;._�nъ֡�q��������:�t�EJ�vuM�(lL��}�e�)J�e��[�LF�tPV~���[D�M>zZnk�ۍK�.De�b8�;U��2`'�v���@�ކ�RL���W6o�V�s��ڵ�茈.�L>D�_��Fl8
sT|d�� �"~fN�����#1�~���	��d�*�Օ�
�蚙�l����Q}n�=r��1<�?j̡���"��(Ζ������G�&�4WPB�U��D�s��h1�;a���Zۻp��u�r�}�fSE��V�Ҋ�#[y��gGM"A����.�d�2����>�)�����|�kx������4"c�k`��q</��`���p737��p�H�@����@�f���X��x����X^�銒�h|��F�9�ȥ�.��'�X����З�}����5��ٴT��r��T:�G8�;����e��enP�Bg�/��0�(���h�ʊ�o�#�7�e�x����\���֞�)�X/[&0�ͷܪ��\5
p�t�,·�<t�o�RU���(RN��ʄ .�O��ݻ��7ߌ}�`9jy�e��3�/ZizX���K�Y�-��[H�x0���M��D$��cc;|�b ����P��HI�Ja���5�g&^�k�a��P�"G=�&��>W.)9 (V�tAf�����N�B�5�����C]��]h;�*�;*�5��!���/o�p֋l�DL�>yГ䬕Jml�䴆�� vln�1H`�����/8w�&��f7�$F ����
�4{z��عs'ҬDT���ٓ6�Cnv���2��&���i���R�Q&rÚ���k&PU55��UEɪ�IR�`:UB���}]4#veZ��<4�!��#D��� �={ɶ���MMP�ۛ�6�}�KcG ��{���WT3�BN�}��c�B?so���L� {���n��*C2�e�a<�=L|��(XB��z���hB~K��λ�(�����W�c�e���"h��?�mz܇��hƙ+���؟� /.�F+%X�|�t�,�P�L*�\'ϙ��Δ��`*��W���{������4�����ҩPz���x������C�VTޥ�"�>�,��4��*��o]��p ���<��>Y��O@^Kr���C�N�v�+��8]���w^窚Z̜u"b�8^y�ui�Q#$�;�@�� ��CS鯀�H ������_���e�4
=�3��c?���Բ��r���f��|�D��#�L*@�
%xUu�FU��+��U�ݗԖd��	�ܸ�p��x"�p"�ڱ\�{�}��k��PO_.X�T���w݉�~�'��_	,���p��}
TV �Ɂ�C��g0d@��g?�3��}����_�
{����Q���ۍ�N|pK�&�����jq�<L��buA�5/���*o�B��!�B��%�y�?g���6���eEQ(���eQ�gP�H NA�b�P�R����t�Nz���@erW)�B9iA�с��������U�Bt�t�1s�����F_�@"�l�5^T���.L�4�d@7�E�]���OfѺ�3��<\�q,��@]�����66��4%��Q&4�a<���Ji�\]i�q�-��oٮdG�G�.�J�2-N������/��	��
�酳�%4[ �U���m-�ʣ��C�{/�ø���2�y�G���on����n���z����Q�!ړޟѮ�r8c�.WJm���1)ە���S��8fq��D��zq��31���%��J'�j��!	�BODcJ¨H&�R;qt*t�k��U����?'�+A1C�!+t�b7�8D���jA�,4ȇ�����.?_ݬ������¶�Pd27
�pހmdB� �|)�=���?o^��Y�a��=I|��r�rUA?����FM<���n�}w�)ʫS���ý���y�<8���9պpv�ݡ�)��c�ǃ��-�Ԩ�i+��}���a E�֩�0���](�5�����E+�}�[-9t,��'���
|\}������>BpQ�]�H�Id���d����R�B�3�`����5si'�����������kB�ʏ�`�%��ɗ����w���7����atn��V�Eqv�j��Z��b+x)L��nWЪbt�[�
d 3-/&(�g�RW]�/}�*�u���u �y�Mؽ��r��o�p5�V��;~?fN��)�-<��!5��UsKҺ(��r�ގ	+"�M��t?�?+��[��m�5*`���g4���Xzp �.:�|4ԎB�>�T�(#S�IZ��Q@������]�1_+U�x��k�SO`���x�V�b��Q����gcg'�)�$,����ڑ&@���6�x����+�ذB����l��B)�e��eT��
HЈ#�U�5��	oKi:����u�4���
*x1��}k�����Ӡ�y�,�a��G��)������V���ͩ?���ʗ�y	˄=��G�� ��CX��4��}�Ql����j��:I?����w�}��3:(wG�L���ƙtx��K��v���-ɣ��2P�Q	 �-c�)����׃Uk�"�Ί9n�I�*��Vg~nRTs'�Έ馔�=0�ć���4�Ǧ��-w��i�J
��%섒�@�sV�3f���.�i�����ޕغc��:��NU5�mI���>m�!aql���̹�}���tdu�)��y��o\��ύ[�ŝ�ޢ�A0���(�6��t25�G;8�$��Ȁ�}�8�<---UW+������7(g���/5�GQ��AZ�R��xȏ���'��h问�$��Ys��#�wŀ�����N�,ݼ������ ��Sz�i��Kژ�B���S؂hTrv�AUe�a=������>�Hl8��_=�����p{w6��Dq��'��������(9���H�S���K�8�ԤA���{�=J:�d�ake3�s�\?�
��Wb�s�}�n����p��S:�g��i�=��(�/�Xp�l��gR\�d��R ׏�m���Jf1����$�}�}�Y�x��M`��    IDATV�ou@`9�ċ���q����~�����-d��P�aa�l ��<������(	7�<�� �~��r#n��o��6��Ig��fF7�ڊ�"�����qX�s�ɪ�����[�@��G]�+��QМs�9�f^#�,QV����TjH����� ��d���c!,s�,E��/�k(`�����pK�y��4�/J����U��\&P-[ŏ7I�0%�cf���g2:�]�$������NDsmX��Tɗ>��cx���$�$r��5�	x���-�JT?���<�k0B#f��-+5^W��;ռ�O&v@'���+��x	�t�o�q�'bтS��v�׬8��2n�8��&`1����8���9�-�W��	��o'_\K>�3o��
�>f���89-t�)
�p�p�EHe^�з�٧�c�8�_]���:�J��K���J0�_6�A�a^v-gR����/������l����7��c���&z��Fw:#��&��:�S�t��������CWHR(;�zp���@T#4�Љ�	D�U��E��h؏	�MO\v�y_��B����Ŝ����ikc>\||g��s\b�AnpH�S18R�w�xY��{:h�C�${v�C��?ؖ������TW_��|�����}ܴ��%k�}��T��	gϟ������U��o\�ק�)og�h1կ��<Č�)*9tbW*��iV�W��墁�|�@qm�j��4u I�E�[~��\��u���a��(fy��N�Q-������`�M3`PN�I����s�e�Aq4U��Ťj��{�wlU�`����~T�][�����R] ���c����b��|���p\y�j��Jln���0y�!��i�� �M��]c�Y+�iG��>�q}�`E�I����7y��c 2�6�9�_un�Τt �
F�, )^�	�3�Q����t.͔I�S�-�.
z��U.����<m@���#4�#��[�<����.�� {¦W����K�($�K:���F���R��b�,9�h@�W�(��\uL�]r�v�6\)��h������JmԶ���V�$�m^�T��/���9;G�T�Fh�[*#�"�VaO�O9^}TE��]x��1�L)���!�Z�i-s]�7���FiȦ��V;#'��}�k��`��F�s����M��dZ�sR	�#����SN���ːg�Ofp��jlF�G�U�l��cǋ�Ö�UPeWM"F#�-[�EH�w����~��4׏��~{�oU@O��45�!���{��
R���fF8&g���;:#!�>��H~�;�O׷��!(�"M �;��?ǁfA�0����+.Z�I�����?����Bgr�e�wf�����':\>#�69��<Y��,���Q��Qh��7�F���:pU��04��`0x����Xu������G�]����h�j�K�EK��vT5����Y�l0��:d�a �o�Q�T�Mf�4���)��/�D���ӗ�sc��ݸ闿ā�#(؈ $�����b��6����ۘ2�QB-=�]�3=�ۨ.�l�TDe����jX���Wm�B���Ͼ`}Cx�ŗ��WQr�D�	�8hl2����&�8}&O����z� ح{>?�V7����b��.�_�^Kv\&��GSC5����~��{�D�LA��3��=��~�F��c` ��b��^��VVa�L�l_j��C�-�+�2�ܭ�����DMu�#Y�e�D��݇U���96G�s��,[��\�R�t�����/Ic;��H��E=�~�����:���)$C�9㌥�J?�L�M���y�UB�S@�ЏEg���Q�j������S�tUK��;
�\���M`+�oS�t�m$���fP卒��\��Ίր2M�%끸'�y}2C�ra��i8u��h��T����@Wo���رc�ET�3p(���,�K����n'��'7�A{׮X��N� J���̀�
z��\�w�Xtι:�:zp��q��C:��r\'�8	/����Ά�9D}%��g	��m̨�6��rI�PD���g>u	��;���B&+� ����׶Q�����݇�'5��p�ޜ䒉 �"���,�k����;�+�M C�OE �@�0�eDCA�k�{���/��w/]�	(���?����<�*��p�\��:,	9"V��TiӉBV�T
6��$&Sb+�3uJ0�hOU��踶+sV-���eK>:TYY������.�ːH?�����O=s����1�p�-\(������M�GP1ϲB��"�h{V%6�S��2xئ���x�C�h&#�.Al�H_���p����v����c���H�JB�˺��*����<���oc��1H��r�������k�d�I~0�[	��_�`����M˹:�vJ��7ΎC*W�����}>�
� D�쎔�{�����	>\���Z���#��!��c 9���`O�BHY�5$]�$��/8}���/!�g �{�?��V=u�[f`0�̘�C< 9�h��U #�.�K+�0�i�g�̄�?��"�_@jXe�s�S����T��R�j.I�h�۲�vP7զi~��eW3���h��4fh�P�� ���c6m[31[����� 2�!���ǘߡ����;��LA����Z� ��&�9��B0ƺu���/Is?�*�	��5�ks���|P����٣�/5M>A�
%�Njh�j��73�q��,�k"år�PXHl��Wb��P�qA}E+�-BeԏH4��k���56ae>~L�֋�
�𷅦l.����0E��DܩL���n�S�:kʄ�Ii�>
�8�a2U(�������`�
?�D$3y�ؽ��?�d��~?�Y�Х�j�}A%�R��Ed���#5>��ˢ$oά)�͏bz@3��h���uصe6��	=ݦ���@2�[:{��<0��r��Hl���ذה�g��b��gG^���
ǐ*{Q$�$^����/�yL�#W,?�k߼b�'�2!�������y˚��u7\������Wc(OҘ��,��4�E�BV��[��pe�ꪂ�̛$-r1sK��e��M��m����Ne]�:��E4�G���ɗ<�ؓw�����Z��Є_��7���"�lA�Q��T�P5��׌��s�6R
SL:|�G�Ă�H�М0����/p����ލ���غc���Q�c��
��dd1~t��{��Թ���%|���Љ!�8;�^f��Є�������̲�p�xH�&4�Q���@�N���g�����C�����ۃH<�T&��&��s��@/"����@��T�!��q�'���}L�0Y��5�ᗷ߇��G��N<�T�hi�K����q�����loC��C�>Үk@���#2��"�#&�ҫ&Q��0E�2tT�3ֱ�К�����x0�2]����j/ۉ��L�F��M��k���T����<��Nu6+{�r��֪�.vD���,�D�-_Qmw4
��o��m+��~-a�f��E�1�Y�o���.>�������=癰���c�),�7`UQ�HC��0G;T�^�����ma�08������XGa�OU��+��)���7��_��"��qM��J٦K��&@a�S����Ng�i�;k��V��RQҭ9�����#��xh�+����*��^xu3�z�%dK�Gg4$����W@��(M��)�faْs��Q��1���>6oقW�xKl����F��o]:����?��íH�Z|��Нn��=�ǌL(��� ߇��#��|/���Ǧ��@�"G�\�����s�%bQL3v�e.���~",�"������)�X��02��'�[��1֛��l��7L�VSc���il��m��|���6�ժ��S���m�U߮ihX,�֧_���G�:�?�L�C��c����}��%Z&���&��Ty��H��"a��Q��t ��@'y�����FT�Dg
9N_���q�Y����?�����-[��DbHfs�ry�����T�����a��&��y�{h��UA�y��o�fD����j�n���B�2ި2Ղ�l$�1R٢�*J��9Y��Rbe�֠]M����Ul2�WEOb_� d
E��r�|�,
�=pg�(���f�kւ����
��_�-Г*�޵��ֻWJ���!_��MI���"����UW�;��:N9q�@_W;z�:��d�	T����V��>L�Ѵ΍ǳ#$B�3Ρ�BG\�4��@� ejߛ�ο��8Jg㕲U��Mht�f�|������n��*��R5o���j��񨭭�� ѐ���=aF	LD)��dD�
�EdP(h�����2i2��o�ܸ�۱}�.̓��L�z�#*7*�q-�W!��~�&Y4�1>���	 &!�GNv�.�I�䜞t/���@V1	���-sVvn�nx��VF�l�Y;�5���x���]�V:_g}}�*Y�_���d����3�|)^�m�q$H��q�;Q��#'6v�2ęQ��z߅��bW]u5�2��z���@�Lp�}���Fb�0�����N���_������w�����v7ti�>y�4%	��]�7�zK����WD���|K]ĝ�ٵ[	#���`b�؝1��T�|�|N��0)T#�P����p~sߔX�ڢa�pv(���n@{�[�4�G7��Ԋ�_����?c8?�l�g}R+��k�u���4l�f�DMf�h:���
��B�R����5�e0g���� �Y�p��D|�6�yvte�E�
G�*+�����~�˕��o����v�C���6���Dp�Yu��r�]8x�hw4`��Q	c��F�WU��*�ʊ���aF͹���vlyw��=����iQ�ҍ����b�g�����[w����?5ҫ�=~Y��1�y~���⸖z�{��|@olj.s]��E��"�ő��զee�Ά�2�p��yz<�U�j��o n>�TB.��:M0x K���A"Q�
����@uM��JbסvQuRi�VU���^dzÝ�C�h|��i�6�׍QU�[�Л,ྵ��m�=��l�;(^; � ���F8�ŕ�_�Y3�"3������B�d3�G|��!�i�$�������g������ʖ�EX���(�8�؄87�ô!M���x8Hb��L��WMN��]q��ʕ������ĉE3ce���.A��H��3ӌA��nW.��uf��pD��\C��<����H���& :����r	9J���$D����B�I�H�}��~�Y#f�	=�=����p�
��M��bG�W�3�<�u���O?�D�C7������E�u 꺪�B�H�?5ҳ�_�i���(%Mg�-V�*FV�κ1	�5�]�_{��,itvvwh�Ν���.A*�Eo�߿
�Z� M�B��1��s�B8�Ò�a/[�����xu�F�s��1�K�|,�pι�a���^��5k��SQ៾�=vu�;oGG��&�|O�Pp0�����ï���<���k��И�h�y�~���!w�SBE���<~L���]x�w�v����?jP�#���*��)�b��r�4E�� �@q�ɘ�ֱj2��r*���X(�#�C���r^K�5	��ʊ 1�R���j��G_�|ݱX�����-������v���։w<�������@(�s�<K4�{V=��{wAwU� ��נetN�:�AxQ��|U
����{��p��_j����0�e��=�%Ҥ���]�`��}��O�}��Q$�k�YQ40�'��q-������V#�*`��{�����#���U��,j�YU]�`$���v����$6�����fEUQU�z��Z������j�լ#��Vt�TF��I�j��������=c&L���O=��+��[6���!DQt邋���"�j��ѿ��'�A�Pw=�(n��^ds%xQX^�{Z&P��c -d0��U�0�AXl3RKߦ����C�2�r���榊g�.��)u�Y���iģ1d�Ic�)]u�0��
�� ��94g����wj�3��{j�
�PԚ�1L�D����y83�:�8���f��V1eS�2>�G��,q�)�ɠJ��4u�A� �)⃝.���URC�mZ����|_|{Ӆ ��t;L���� %�4��%���`l�31ȳ�chM��k&h\�bY/g"������e+���I"��w��k�����A����Y#'�be=\��o���9�l��7ߣ��{B�V�L����b߅#G�����QSU��˗�q�Xq��x{�<�8�R�yQ�%��	�Pr�A�2Y�R�?��՟�4.8�~�x@~�<;B%֥�n4���+����[���M�2�?��ߢ�p�����j**��^z���V��������t�x~r�q�9Xg�}V�\J3KՏ�,G/�LL9��Խ>섊��X(���x��3���/^uL�<�����%��S��J��ryo0�Ulҭ�	�ff�l�x��Jf��(��Kڸl�2�+Ѝ1�D@J�������?�%JV6������#��FUߞH$z?�\��)w�_{��Ξ94X4�IM�~����x'�saLu5�O��Z�����NreMx\�3���%	_Z;����a��6@3F�����u�_�3�8�v���~�3�uv�*���h^�%d0@�Z���o�M�����z�}��i�9��98���
D~ 5��D"ر�}���ftvucڴi������3<���[��]K�V���A�Q��XR��--�v��Ȕ\x���}�$!���i'�B}]5�|e�l��o��Tw�ԍ���V����*�1��?��?�yl#�Ҹ�5�������G���<���`/�Her��/fR��LU.G[���1ԩ��*5JJ�$�+9���
�H�+#54�Ì{��5C!��niӜ�l���řa���Y�.�[	y�D��(��� �UK�A�	���e:^�Τ`n˚:�.'�u�V8f�b��
"���v.-�1�nͿ�E��|�غ �jTUj�~fN����C�z��n�k�ܩ�Xȫ 	Y��C���ۃ��J�W������]��d=��>������DW^q)FU�T�Sw�ƍ�1�e��"�5r���I�������v����t��2�qP;�:��sY��%���s�ۉ�BA��t����l~yW E&��!؝�&�^�����Ԓ8��yxx�j<��3��1�PD���ⲫ��Ɨ7	�j�yv�:¿���w��\����k8��LW�N��`��
i�***�v���Y#)n��Q������a���Ad'��I���-�����y�Q���'�rBSӮ�O>�`Y�<[�L	z<�@0X�ZV�*��V.�+���b�X�M�>�<�޽��u��E+�J}��3��Z�g�.�\���G=�?��Yl?q�RNVy,��/�c	�VnhZ6���T,��M!*oj���.}b,�����J�$�D� �B���V�g�l`����v<�����ʊR+e��x�#�؏��wFkk�|�k����&ݾz�m;w���BXr�B����;nE��E��FCES�1���<�e�C��B��A�:�VQV��fИ��7��}�r�z͛��Vkӄ믿'�|v�ދ��t���!M���-n�'	$b��!��6�÷��k476��Oc�wc���9��8g��X�h�(f�n_(���lݶ���SK�������k����Z6�Ndu�IŬ����v�̖�$K�_��N��]k����׍E���-S�1�*�J_��6�<���F����b��C(2�����?�L�<�I�v�Z�v�j�(Qz�&0pc0�ٳ%!����N��8L�e�����b3�b焭qU�ܞe�*%uǌ�X@�&6L�x����T�FMO��~#d9�x���}��,���S9ҿG%������,�"V��x���垔g    IDAT�
�z'&��}��K#�@��JE�)�>��;q �����w@iU��>{��O/��������b�-5����5�$�H,�nb�4*�b�X@�Bg���a�a�������y��G�����s�]�k�`������۞B���]RE��y�W.\>�W�vn��iJ�<��$~	�\��yNN��-�A6�D2�dM�����^R��z)tw��C��T�=>��Z�n��vД���S���5�ׯ�_|!v�L������"缜`��^��3������:΋�_:�6�˩ڥ��5��$�Y�Ι(��}�GcԨQ�۲u��*�[a��0�0u7x�a�!���Jv$tw�a8�����҄�[���a�[h��������"�J�kЯ��2�����桷�K�:�3Ύ������Ҧ���jdQ������ĉ�����(E%��b�hkE��K�q.��8&��3U�����;ef:��?��Q�m3t^	��>.����l��U�������m�uWg�0V����y2��̮D0��4�24�+�v�Ҧ�$���%�.�	k�@���i��`�i���뜅V@T�LC3�O�д��mY���c]k��k.�Kgvm�0�r�\.��i:Bb�&|,�ïi�ç�t�<���Y�4[��pm����K4��&�gzF���M#�P�ġ����Y+{�t��I�U<"�6sF���9{"���-"J�pp�qDҎ���OVdv���=�G"�{�**)))i��}·k�=����l<,�ḣ�Fee9y�a�)�aY�3Ę!1��RZ�F*.��h �hȇ��x�n�������93w�B������O���Y�H$�^�y��1��ЀY<�u[�"�7�	ѴFɰ���b��5�<W^r1���f����Ob��/HK��RGuN=�DT�W�As	���@sS�|�����\��x�u{�W�Q1X1�e�Ͳm�\��N�G�%������� �w@����v��5�p1]����pz0�؇P.!}ܘ�5�>�X��LjF��3n�����ځg�/�3���0ui�"1���yaEps��,���=�"�KOm�e�
J({l'sL�6u����%�L�R���&�~8㤃��iS�J&`���ր�n��17x-���R���7��lEyc%$�A��w����,�∞��	Z�m����E�[���6�rv	i9w8]�U8�v�Qos��Ə���" �(�?�uX�s3O��QQ�:i��'�S��p,U2����Y���}�Q����B��X��lؼ	o@u&^B����n� ���Z���X'$V�P�X��.{m-��I'���8�պ��Z%��G���RE�:��	����r翥�u{D��Qi���c̘18ᤓ��&��h�j,\�zҔ�l��v&�x�!- G�"�n��l�%1���q��	"+��6���Һ�~�%�|o��[����׀�/8F.�������c����}G֍m$r��,�뗊���P+��|0�M�&	�I���8Z�L4�ס�ez;;��ա �������񹴠����.�si�����VӴ[�����q:K��ϭ���SG���*W�u�ʟ\�F;&EѴ��v3Kp
��i	ZT:h.���2��k$ ,���0E��%5���tR~[����d��f!N�xڹU�a�[�fY���
��ʦdȧ��T:����"��k5��O=��!�����5����]�p��D��b�hZV�:hv��)d),b��]Vfuٴ2;ɑ;M�6<+xի��P#�	��v�d�F�	7BM�n������G***�|Ӏ���#�=��-�MG�TTb�ԩ�����O=�D�K*�~6h ��J%�R���$�'{;QH%p���<��Tz�n����`�^��/��PI� ���/�cƏAs�n��������^d5*n)�*�y,��0z� ��������ü��Jk<�u����9g�)Jn�
������r��Z477��w��ʕK���թ��p ���"�v�Ft��a��&��8&d�%�菋~y)�k�=��K?B��`��}`y#h��������FU�#�t_{��Q�(�s�[n�#�?
-�]x�ٹ�3�$�
|��iHAg>Ѹ6��g��l�wɺ�O��'�3��m�/��d,�D���-�!�B7�BAy���eB�dk����q����d�1���r���t�����l�Ma�׎0������W{{;֬Y#Aݮ �>��%sx;��9�T"�}6k�`$���dN���͖I�x>��%Sq	�S'O��~v�h
�����������9kW�B��Cy׉��k�I��H�G0����c9{w���X��g�硇����PL�dQ0�g2e�RR�F\:<���XC�Ǐ�;�L�J˱y�,�}�{�d��900q� ۾Va�"�<��Qb��D�M@�J�Xe��lI9M�S"�*� ˒�E��A8��cPʄ��k6n�K�.Ķ�f��k�5���D�#^C&��R(&��v{1j�PĸoZ�q�̼�W>߸��V�Sq�|^Kkg�ｽH@�<n�p B@����f7��*�Hd�2h3	U�zX<S�L��'�ܗ����E�)�Dw'v6ԣqg��x��M>�E�砤���˨�@y�l>�0��0Ѳ��b�ʄ
 �^
߰�PS_ ��G8���}��{[X'Ipl&��O�õ�"�'��ѕ�ja�(�3>��1Gw_k�!8�=/Y ��t���"���x?<t�o�N���7�S�M@O��շݞ��8�	讒�H���� � �tf��*]f�4��gs�E�p��#\�p6G.:�q�����/�Q��4
�ኃꗇ�����N�t�����K���k��<A�����຺���,YzӮ����EE�!#F!	bK�F�8 ��f��O'���@�s6�,u�s���P�e��I��轇����,��Rx��̙��2d���
�5jv45J@����&Le@�]�]Fc�µ���+�9�y�̟�����^N?�d��9�Jd��ʍ�b��TU�ټa� v��}���c��w_�#A��h9��3J� �W�Z�)L�
����H�?�կPZ�)X��3���E��
��r���*�r[��0Ni($]�]�[ehji�̙�cʤ�hj��3������"����H�2�\�¡�ɔ��hn�.����~��f%���J�Pn�lZP��D��{B���YQB��`8x`\p�y���Bg'��������0P+����>��T���P�� �Ug�&�kn<T=#0������R�%y�dS�͈ϋ%,�	��YPm�B^��ec�j�N=n�4	zs>��W֣'w,�8�I�򩌈��u�����-�3&�aQc��X�G�rҕ;��<�IN��Pk7l�]�=�-t�=]�ٲ)2k�e�"uR,8D=>��>}F�!A���������JB��B�Cږ�jw��8����,&/��i��O&��)�RbF8�'x�����Gtx�z�	iS�|�i(��',�@8�����>]��ޔ ��=� ��7�=A�#����%y��teq	��7F�X($����.��>���^��]I��P�-��A����~z6<���^~I��4��1h��;�@�U�ܟ�=:σ�6�f�>u�T��}�+<e$HĻ���;���)׃�9�pBe��L�B�y�$�я�-!A����^���S%�6Ŗ��_m����8].�F��ęS)eAIHm�c����c�+�]�3�;�t�����H���:���=5�sb/ğuk���\��O����&�wuun�t3R����u|ЊBpEB��;�,`�&��5���`��L�2J E��	դ��~��B��E�7�d��MZm��Ղ�,�쉘�K�J�)*-��p�d����*J�-�Ǔ��rnò����Q��r��K�t�h�IE�;{���\ii����*Q�_͓��qC��njZI+���eW:;Z����\*��m[�=q�X���*�H��ԑ�==����R*�*q���b؈��7�{�z�nF\g��]$����Cpݕ�c@Y� e�{�I�0�9x=n�M?��p��	��'�%�\�R.嗼f�:	 }�駂�6|�,Y�SO=E8�V?9�'X��475a���,�/� ���W\�Hq9�9+�X����0\��+��J����Q󣚊XL:�n̛�6�n�TR���L�v �ۻ����xf�K(h~���Ո'�R!��F��I��[I����W-9i/����|6%�o�`�?��{)-p��H0�X4"mP�
C� Ǝ���
�%���;%\����HeS���r6P~����i�:��ٝ�:+h~�SI9�y�L^3Y���Կ����M0�I%d7�];`92��z'B��{V�ٌ y�g�y~��|���ADJЩ5о�U*�P,*ɂ�pc�u�\V���@6��{���qD��{�	O ��_�ŝ��/���@�:!A�"����N^as ~K���c���i``�j	轝�ݸu۶���CF�HP�3i�
��*v�;ǾU]w��M���O^g�`,$k%�JP�|y��Я� ��d�3oP:��֬����
u��4����+�/lASg�`g�+�-9�LNJA�r��8��K$��Q�y>|.���_;w�E'Q����%���bޜ�����R�#�6j���K���^�N�Й ��I�e�QGɵqdp��D�����Q_�=�]��9��N����3Rb V�{���-S�>��=��Mry�aE�����}�ם�쟓ɞ*�{|�Dё�0�^P|K2?��(>*M<U�����S_��i�9�<�/��c{����t��#��7p�ߌ�g����z[[�iÚk����z!�v<p�B�Ƣp�ª�p���M	F�2R0��5�OI�!*4� md�y���y*��N�7-��!�}	��)�#��������(�a�a�2����,²,�e*��C��eOIR^�ggWo� ��P$6Y����p�HDd+������CMn��a.�g������hC2�#3]Vzu۶b�1�p��ɂ��4l�ۉ{y=����j���]�{�MM�1���ہ�N�dry]����:��.(`��!���W``e9
���!�B�s�p�9g�ܳ"�T?� ��%���:s��߿��m۶aٲeX�bF�!V����.��}�6�]��.�/�A*'�pv��ፅ����k�G���ك��})�To(�Pq��ˠS4ۋ�υ�̺sB�z~�|�n��ъ��p���`ځ�E��R�?�,���a�-t2	��&%��e!��9��l(v��U�u��K�7f�b`�fR�M���U ���)��L�-Ev���T�C1��������l(N{өȝ��ܔ����'��~~-���Z�Lj�Zg�)��W�rε����K!>o����00��l��AQ9��)���>\��}�iiɜ_��8���8�����"Gl7w���iI2���ݠ��������[�l؄{xuMͰ�~؞��|l�ӷ^�"%�<����D|��`~ȡpY	|L�֮]��u���	� ���Gu�B}�!a���g뜇�<��DbR!�Q��M��A��L&QZQ�	�M��I�#��".B{w/��=u�MHK$�އ�����B $�(�|zy3� .���U��;jk���w��ܬ�ؚ)��G��>�&�X�k�-D>��^ȡ8��W^.	��/�CcC��BP&�k��`��u�JY�/g���1��y��-�#�8���lH�L��۶[����MH�Ta%tJVߺ=�)h����s�.�׭���]���rӲ"ܒ��2��(ύ�)���k�I�FRQd��̂�h+�Q���Q弝�qM�voX����ENȲ4�n��?Km�L�-��!(�/��˙˺�1�F�����LK3��0�����M�Q��>~��t�"&�$n�S�x<��4m[���5��6iR����nm�׾��l{���| !ZQ�`I	�pHf��t^�E��Nu��p$c�H}(x���2��R	"!p��N��Hđ���Y����v+�j�nq��f�.�W�&�����j��`@��\Ф�$��t[G�Y0̀7��'V�̲	^#���h��Q��dE����3Y�ti�ɶ)6?�~�;��Iĳ>�b���
\�:{�{�X\u͕6|8�66��Y�`��z���{E��C�=
�p^o9�?���ү
f&�g�|���0�g��T�t�qp�榛��yd�E�r�9o�X��;w�a���Ǎ:ۼ�sp�`͚/�a������&��>������QYV��/�C�GK[V~���qTT� �JK^(f9�"�Zs��R<��|��|�Le*��p�UWb����d1g�x��9Х�ld����)�J���(Y�$��f�S*sN{���H�K��Zpʿ��4@�[k7���U6� �Fv�	i?;��÷v@q�N�vP�N�v��#z�*�T]�=��Q�r���MQ%�ZQM�oW��т��6:���2�ǊJ�y�Z�����*��j� 2/h�c�U@?묳�ڽ�`fΜ���)AJ�`�������RĊ�����]�TF>�6͍ϙ�&&O��[o�Y�/�o�]�>��uBCd�/�>�W2���#�jf�.>�>3���(��0�F��uDPc>��Ν��ݲA�k��4>>V�|�C������Z�1�UCuJAm+��d2%�C�1��s�߀	xeUUEcbm���	o���lCGOBU䚎4��4�;^�Е���N�d��Z����ǩ'���|�^})��ؼ~&o�G�˯�kw����Q%���Jqݕ���>w�shiޥ:%�r�L��d��t�QG��k��8����5��ѣG��0��j�nd*����$���q ŕ��(5K&L V>�;I�G�iKYI��~��]���\�R�0�LM�knWZ7��t3�r�!��b@d����偙�iB'��a.]�X:e�]Y未�g`64��HD-�U���mr� U��S���z.M�cZ�W�,��[^����4S���[]����B;���l�x��\�e�5���4���-]�
�����)���E�<��i�5)���ΓY���w|���H��8JE�R��c�]L��Q��7]��ek�++"��\ �A� r�i��A�5EʤR�����ġO��p����! ���Y���8�c�ˡ��¦%�'@����YK����T6/ �ްr��%:9y�tw�jA�$��
���SX�* ��C����ՓD^���g����ې���F���������:�u�=��ԂY4���H4")�8���_~9���|&�'y�����Y�1�y���H�I'���h��u�#�L���D�m�[[Ű�}�!B]Y���r�)شq=6�nŏO?o��6��=6lF���='�_]�K�؆���5���*��%e(.+U ���P�	�Ҋj<��l��b���T��n��&M@GG7{�,xm�:/\����G�A�;
M9@4�彳a��l�̟	�#���7u�)CJ#��pHd\I1�qr���q9;|o�;hmU�b^?Q	3r2Gf@T�?U�;�׃�׳m'��d�:�l~��w��
���2W�t҉"��v�2>���F��J(���ji�s��������e���C��`�F���&�!I �;�<�0Hϟ;O>��T�b"�*U*tVn�8��&�-LΛτбT��-M�2�9�&��WZ��V�������)�PҞh�bk8��r쎘� ޽�4�^e�%�<iF���%ݙt�ͻ����(�<��#��׆#=A������ad��g����`]B���`����INEh�`J���%x����p�pyarv*���X��
�J�RUb�N�
n�;e����K0���x�������L8) +-����흽�5k���$V��ƺki    IDAT�A!��SO>���-v��8�\�*!T��3fp��JJX11
";���9�~:3�qE���0u�)��n���p{�#½��b��S�E��0v�_'��;---���~���d�q��`�d�=�h�x�jkk�N;�4�&�/��������2?��ϟ�-)/�x,~zS�/��Db�r�ܩ�}>�3b���wwk	�ߘ4i����;��,�7��h����(�O,�C4D J�J@n4W�x!S���V� 3zn�lAx���Fa�H�L�L1D�$s7���%�b�*���:�p8*R�\������V5;:[�%��`�k7u>L+g�i�f�Ե<�5t�O��B݉d�^
g��ЙL��'"화���'<�|2e�E�R�1�	���
PT$��	�;�Ů�<����Í�x�pC�ÕW_%}�:�y�}�ڼ&y� j�;*9�YDH�)nk�]y������?| o�����p�Y?��M��Ŷr�7)*t|�8k�I���{K��شo��>����k$ƌ��^Y�����=��x�RL=`�$-�<,~�-��A���KQSS-�F&��sC �f��A��z���Jm;�W��^Ɗ/7HW�����G��C?���,�,d�(��M�䓎ǉ�����,�Q:hmm��ի��G(FSK�m���u���1h`�Ċ$�`�~��e�s$S�Z�HDsTe��	��^8U�C��U�ܿߨGOh1�"��42p����.�g[S��s�=U˘���<b�0Y/\�<.�f��S������2��q#�ҁ����	tg�n�4S�V�9��Q�Y���9�\	�D�ϟ3�?��|._�\���9д�����R��+�s���A[�n�fwL|�X���0v�h�}�_%�X�~f��0�ַ�Щ�ǖ;Uveg(1���\^݂���Y:GY�%�؇ �CEA.@����v4�ډ�����	��	��CaA�;ʓ?��(PC�
(lII��4:��("E1��B�l�р�?X��+>AO��`���!=V�uO��̈U+�(pZ�[7�Tɥ���p��b�����d|ǟ����lŊ�p�?��{�W�#���EE�y���4<��3ؾ}R��4G��7.�O��T$�ǒ{R��N�%פ��V��bj8�K%�2n�cKY^� ��W  ��53����aH�߯���çM������]�e��"��?�/W�;�W��z��Y�D��"��W�@�
��y���HQmDf��P�U*�3�ϋ4�z�1�^tf�HqH.?ò�I`��-RaWWWJ���aiq�-?�����˰^�'����B>gX���d4M��|�P X�y}I��N�������Ƴ�h:��o����k�I�ҥ��)�Zp����+���ʜII$Dy,��`%� ��� ��!ԓX$ �n�����!v�w�E��źMpB�.�M|�ޣp��cȰ��khĝ�ރ��M�{٭���b"^�������+~��������x�{��{�J׀��Yg��)S&���L����7���A6�4G0������Ak[^|�e|���(��d�ֲk�Tt����6m�EGO7F�5�&���g�v��44���m;���*���£����M�X���J�Ĝ���k+Яf .��
8@�C�����&.n�9����QbG�&��H��$���~�J����]�m�6x���%�J��"]�^4�!����ŋeM:U3AQ�9�+�P eG��b$���ȿН����P�\�W�kڑ^��u�/�E�Due)�;�XIH::;%a�ޥ8��ot��qsu�I'���}\�� �&��.46�BW<�O>	^x�����<��#�<MK��|
]�aܸ�1jo��J���*����Vn���(mtyO�o��&������w���ݴM�� ��������J��@"
�\Y
Ͱϩ�%ly4�}ǎ���#�+�>������CX
l��tL�Ȋ���X]��:BZ�<w�cr�y�t�olƊU���U_ Y�XPG�ֱ��Iׄ�"^�rfNa ��)}v�X��f!�?���8�Ѓ�M�ѺK���1�tO�<�Yُ>��=����+����?� bJsf?#,��}��?:?��1�	�r�݉\�}j{v�� *�-moUC�&�"I�Ig>?�K��!㸂��ՕU��=쐋o�䂥���o�
|g��X;�S���������@��*��mn�RBiDA��NXU�uG���pHq�@	�����(��@YU��T��,V}�
��<t
q��Voiii�K����O��v��Jh~oҫ{zM�0�:
>���x
���Y(T[�w�(��C�0�V���lon.�r��ɋ��wm����D&L��`����Rԝ�,��>��è**�j�2Ei8��[��h$$��H,��t[wucѻK�~�VQ��>�|<�\{5��m[q�=��ng3,z&ۚ�4�җ:��fa���7�����Cp�=��޻��[ ���G�C�.2�-�ͨ�Z'�0�I ����!?<�L��B[�R�M�"�@	OJ��V���W�k9�->��1�L�2E���>��c���"��^Ç�\��=�M��5���!D�*p���kd�1p�`\~��Կ��A���G�����1�)7�yu�~�Q�77�e�vq�"�_��G:!�����ͧ��]q�=n�C��5��$Ǘc0��k�/�;�T�ܠ�>p�c4���sg���7�j���I�d�c�p*z%����N���*.�H��N�?�Y�֓�t	l"]�`'��9JP`8O�I>f�{�[�D�N:g�u�t�-Z$	��i	��ǧ�.I�l�W���-uy����wuK"FJGG�z{���F���w��D�����-3��v�hsM,����9&O�\�QĈ�P&%����f���8���1z�Q2~���fL|��f%��Y
�V'^��P��!M�	�Ǉ`$���$�U��h�=�&�d�t������e���W����by���gG��>v>Thr=
�^���f���8`�>���I()�٦'
�����:�7�d�R���;p�J]�C��-	��۷#�I���r�'�*l��˨�/�8��a~}$�W����-`D?��H��\����b��+�����1��n��yߘs����>�;��U˪׼���`.RV��Q�F�����%Ȋ]fIv�ʇ �, f���
�3����(��@%�M- ��a۶�qSa�΍+������ҿ�J"_VVk��ھ쏾����]rWCc��hQ)~0y�<��zi�
�|//�a��A?jJK$���M���X!��H��زc'�\���:�t��

�/n*��\y͕0h ��m�̻�B}S����!
��]�]f��7~͕�.-A���x�A���"�p�9��i8�����SW�����֊�ݻ1a����e���KlݺUtTۙ��
b|�L��ٱ]�j�F�����l���6m�(�/B�s���c`8������{�ǧ�7�t�$`�����a.|��ǰd��Ȼ��z/���� �]�����ʋ"p�\^��X+AeU��� ����d$����fr��͒��>򯽶���� �����\�m-�?�+Ou�rw���{��v+�g^��3�r,��w��Sqc8��s��л:;���s�lk�vii�$Q�,�th&����_�e��i �bӖ�x�ɧQ[�MLR�>�8㬳侾��k��p��k�M�h�b̀b�O&%�PI��\��%���S�`���"D-���Jʊ�Y��3�qK,�W�dk'2�pkF�|2��P�� =�W�%P]:��!�G0f�0b�`�2���i1�!��IN٤�v4�M�]�P��C\�&zz"��{����iܵ��_�߈T�@F�ч,t��2F�EǜHo~�`t��.|g1�QI2'ڢF�J��aQ$ Y]ΨgO!�(H�i'b�)������;��z������/e����N�MQ�s��}b�j�������
~��q.�T�d�Pd�C�TPO �4m�G@�S�G����ACꎜ~�������������3�N:O�~���:��n�R�����b���C��HeR2g@���p��А" �뇷�H{[2���-������\6�����z$e�g��!8p�Y0��>�������Jj�}c�W��9����y���v��O��aڴ�$X��֛,�����6(LB���A�4*���ij�E�@�];w7�v[Z:���)~��vy��		�������� l�߁�n�M�ۑg'�(�lF�/��)&1y�x���ע4F��=p�p��}������/���H���M�dn�͚�?Q���mG�Th$�M� #5oS�*�����S����R�϶>�H�J��?���J˰�>�`��&H5��4�~a���!C�������0i���|�'���������P}8h�~ܯ�+���LIp�K��d���|���f�|ح���AU��3��U��觟�@mm�lxk׮�;�ߒ��qr�FC�5��U8g�k���:��s�T[�(����ug��l�{&<~��Pm
��1r���d|�w����W]�Oպrɸ�1��WS#U:�T�͟���!�+�H�4���=W���_ģ�>*��2�^z)2�<��[-*��c��A��xO�`Ex��m�Ub��� >]�����63o�E����F���;���T��38Ɍ ���`Q�����g�H�`@�8��X�O�נ	����#�c@���BI4" L�]�N�әn�ư�!
�<��czI�'�7��U_/��l�BW<%fEL�]���Kd�+�!� �Jث�|�j��-�v�B��}�D ''��2s:����Ҵ*�-ubw|l�r�_Q�Yw܎H ��_{Y���m��h�k���ۇt��[ۯ$S�8�{�4�Zs���5�[ �*&�	�"e�yH���~$H����)Ϯ�۔�6hp��xޭ�<��
�[���n�Z�ݴ�xK���[��Fp�ǤA3T���jV.Zo�Tb�Uz ���$g~����%�Y1qa;�?[^Y����u]���_:j�5����������䃇����GcE8蠃�޶��!Y>�Cl�+S�����~��p�/3�T>�L���z�.@W4'α)j"�	���W_-�i�w܉�������X�&��y(	��x�x�5(�2X.���˗,U<cR�tR���w�Q�޵�<Ҕ ����P� [��M����\Z���m�*�7�U�Y4���R�ũ2��}^E���'� �L:+ݦ��r������e��~����K�߾���ю'�~��ǹ�n�A��h #�����$���x�	��t&/k�1�)���@6��xw����n�رc��]�trye��f�NŬ�y���
���+��Ӫ�d�ϗ3�t*lg#�u����e÷�ڬ���/�N��lmo&�ހOT��\?�3���S��˵����g����{�����%KQ��Q�;+���;N(�<����㩧��4�ᨑ#qÍ7b�ز�5���豣����\��	$9?��?�0V|�J�#�8���FD�c�Z߄?��l�k �zt��gUb�����L�h�� 	�5QL3�U�iH���K�qV�4�2��z�HEᐤ�?ҫ��S�ƀw�[�A:Z;;д�Y@�������Ѡ��U~���ǅ��S�ױ�U`@%ZD��AD�t�ĕ���m+��/X	�Y	� _A$�	�#.FP9��`v���?�4Ë/�~8��2������ѷFU�Uk���:��3��?U�
W��w�Ǐ�?(�����;�G��F� hA�](t��8���iSΞ�s>�6���?�N��_\kժ����O�in�,����/+unZJ��"���8�aΑI[�Q���A�T-��:�H��(K��,M�������=޷"E�wk���/W������Ec�\���]=��B�"�\�;;��+/
G�؈Hn* �p�O��b)�&v�Os��?�L�\[�<d�P���nE~�T;_|��B�h��_���(�
�l^�J�8{����CTh;	������;}��)��m@@MR!��+�8r6%�NIX��������a�Fu��Y���,%Y����T\͔�	[�D�I��0n��P@P�i:�y��M�x�#����LFuy��՞�=s_y�&g�.д�(w"���"�y���$՜Y���9A�2A�1�3��C�W�SC�Vc�v�	(++-{�сA#�5����E��v��p�?N��?����8��":T&ӗ�x��������t��U�-�!�[�V�B�r��^31������g2̯��&I��.�!e��O:�\x�r\/̛#���ơ�����w�-��W`����'b��jd8]�k>���YKK+:�z��3�c��M�*��i�0�?"cS]#�8c�oێ����.�P24He�O�[᤺�< d��̒bA3ho۫ĥLd��c�}�))��h�PX:[5��DE��;ԝ -�
�̹��������6�V��cm(``{g���c�b	�d�2ߦ�`�l$��噠�ν����)ZL��nQ�-o��D���Q!���$&��O*��pӍ��^C���/��*j�#�y����Hg��C��(�N����0
���?�aW{:SY>R�������"&�9��?tڔsf^���ی��y�����H]�΃���EF*��V0�C� y{2��beEI��d�T�"���2����(�Hy773�F��a��P�K�4����ť�蚊�c�c���yk��/��\gw��h��s<�:��բ�T��e�p|ʇ���{�4��!�C2Y
~�K�b�J�AX̠�j�ץ��J�\|�06l܄;�v�辧i<B�)��0�憐��,`���?�	�a?:�{]�v���\�zU�V��������ц�ݭ0�҉���i�Be�u[֬_�~��*Pe�bta�1h� r�4TV������f&ϟ!�(RT,�G!��3�
���Ѥ�Н��A*���HYIHf�m�����7�BJ���	o�ʥE�#�ѐ��P���CNP�}�b���"ҡ`F��L<)Ւ�OV)��;i�D���.^�vi��WV5��u6j���I:Վt/l�jG��9�v���$���?+�E��]��g���ٌy^*�P�)�W�dR#�J�t0�+e���L�:� Q�e8�s��/�gh����'�d�����˯�����m�*��?�я0p�x��X���F�y��Y�˖�Eo����n���I�샛��Vjm}#�t���P�	����(wb5Ri�ް՟7�ho�.�u�9�4��#�	X��UR�\��/74S�b�b"�C��hVx=H�3�N5�s�th�[�X��zn�$o��C%?䞳ÒW-mI�u�$����3�2�t�7��募��2��Fmw��y_��'֠
�!�q&��سY1��Ӑ1�bP,|u��ٍ���+0a�X,~{���2g'�]�-lʥ8�Q$ɖ,���Ka����k��Y��I�5,�'#��@]�v$Ӥ�v!�B��G0"���,���a�8r��so�>�k1J�ͷ�i���@�����:��S����іaVQĤg-�BAY��C��ۏ��	U+A���c�3��{�u�{��k�5��#�?�����1���8������y�f���q�w�	'c@E9�șא��'����!R5H���ݐr4��e\@ꞃ�w QX
�"�q�f%hP�'�}��~�]qQ^"�S*�|^���o?�gn����*G*��^��)�	�n�T�� ����R���� �)ө�r�o��� b����tfϝ+�����(C�V����$����F<��wJ�DjR� &�) �,GJ�R��0U������E�]Vh!�W2��������r��C�7�+�tCf陞n��M�J�5�)��L9�x��@4���=G��͏z�?F��h4�OV�Tջ��dYG�U�Q;9R��w9V    IDAT[�N��|����e$�V "g��ϝ`���9��?���S��e�$�)FD*��v4��nX��]���(Ԣ�gV�"*b���L�U��$v��g�.�u��������Fj���0����D���Ɓ��3ޡ�z4���e+���a�V�~�&��?^q���jw���3����F1�!>F���T<�~���q�����6ږf2b�����F�ګ��/	"�RY*���t	����z��5y3ɔ��S;a��2of�H���8�a ��8tA�:x��b++��@;w���	N��R0!?�_{���4���h##
V��WmV۔7e�,�@�!�9���݀��!��[�+i:l���ڲ	�W����?�`�x�Qi�;�LDyoED�O�S�`R�|�\�N@���S/�8#�텥K��~�N�i�Mp )\g�X�.�>�a��!��5}�y3/����������j}�_&��/��M��k��P��-+����>�O79|r{,
�5��+דN't���`b�'�Ye���vG�~�رc���w�z~Ŋ�G��7�7�=���?:�P${���avK��3���n	�n�E��F47�k~��rii�;��\F�>E��HV
u�>]�{�i��`�b$��s�"F�_\�34>�[�7�]�:)���P6�^�p�HeҢrǪ�t@�Y�!+_��U��윹h��}�ə�+�s���ƍ�e��T�ש��V>h��fG��	���I�����B��h4�񅔁�aJ�5�����xT!�}ai���V#���+Qd�׃�iv2
t#W�3�<?,3�W���` �L��#4�5;f���.y�}	,<V���8	�c��i���+_������i_:6QM��;�&Q|	�7�)�78,�U�Npw�3j����v%�=��F�"X�ʙ�/&"}�e�Uѵ�t����I'����?_�U^z�<���e}8�KS� R�O�)X�*]t�9>���H�#dٲ���yH����I�r�0fn��j�E�q��4c&�5�G�/�ݧ��)N?�d\t�y().B*���hQ�=���C>�o��e�A� �,]�~H@|��rW����������G#�����
�����e�5>����_�J����^I�܈�x��'`w뭷b��!ؽ�U,l)��s�g_`�]��eᘗdi���2R�왎JsQ�P:g�T�LpH��$���i��& �A�+~�+L�w<6����f��X����b�ҍ��ջ��pp"����}������l��J�ˠ��g�}�Ɲ�DL'^��r���Q��;�1�'P��P��eݑӧ���\���[�Y�-}���Y����*��\�2��B�Pd���uh���<V^3��e
��]���gz���ݷ���о�����UՏ�e^c[�4΁G�Ԡ,�'��n�|��8��)eI�>7<:����:i?�]$ܘ��7�ٌ])20xt��p&���Z�w՜�f
�JW^��2����A�0a�(���lL���A��)�n�B��'�!�<�Π��lJ@�4�����k���=�B��Ri�
"&�@4rh��CX�`���#ʹ��&*"��v���v0{�߳�A�
�2����j�DC�n$҆8�I�^����^X}gRqIX�R3z"����Ӥ|+Ĕޥ�mO�n��	i������L;p�(�-z�M�Jƺ<Ν�r��f��g�p*wg3t6A�؁���8��k������T�N{��P�*��}�>A�l��g���ܪ�.��-��n��� %�,2�:U�r��H�=V�r�lg�y.8�g�eNS��~/evC���у�(���jt�a�ҙ�$����09 �|������U��>cF���]+3��;q����"���r�yA�ϼ�V��v���d�x�y���W�G�x�|�B�����y��k���Ï�9������AC$i:cQ���Y�|�����uKI� mp�9i-Ϻ�nTT��G����-ҝ:��31�����c�(.��"����!�#�3?��"ttw�Ιwb��+E?�`>���JT� ����q��)�,��<�(��t�(���h���`�&����	l�v H!��I�!�L�%���ו�x��{����("ZJ��1a���d��74�f=��o &�)}k'��'�Dܿ����{��~�M��������˲�wc}���fI� 0��ԴCU��oz=�����^}y^}[�Al[��.x��p���9f��z%K'%O��]:��0�L�&����n݂����K?xҡ�&�U2`��l�4.f粑��Hg���<��D�3�O&zEq��z��1�3�/�ғ�)�C"���m)z��ED��`��~^����>yP�`D���&z���(�]]B�#���>���A��@![�����n+��~����c"aӲ�IH�)
[nēd��&І6
l�Ԃ3E~��t��0nX�H�F��J[���X�T�k*�s{
��$*�	-8���)�蓕��n��Wmj�t�{˖�Z�N�b�gx\�,����Н��zn����Þ�cg�)ɀ�v5E���I�1�)�����J��<���x_����ű�[p��u \@��u������z��[��:|�>�BA�D����m	D�D��H�-%IEI��H��
J�
}���q�f��1�1|(n��*�mܶw�G�T*!r�d����"o����i'��V4l�!6��ӟ0��Ixv�|���JT*�7���j�a ߺmn��v����8����\�˟�SN���?��s�J�ˀ
�:���ˤ$�S~���@Ss;������ �X�������ŗ^F:����)���ɧ�A�`���?~�QyNn���yK�<�lY�w0�`7��M�YdEQ2�N��8��`5*�ql"�?)vAR�C�U��R4���^��{��'-ǒw���Q�U�z��z�=��S���~��0@�*l�G����jp�SRQ)4H�-����"�p�V�]��0�%�v��	(��!5��5}�9��o7�������}{�����ym�܎�9��bW.	3�#�-�O��ɽQ
�K*t��=�t�q8���}�Y,\�y���4�����+�P���:A.�Gٲ���T����4��Y5e�qA���N��!�P��\9@(S��8��VD,���[H��Ec��Yt�3-tg��oi�'k7�WT�iz9KW��|]CI8�N�������_���1[�ܐ8D[�� Ќ*t�K�T�T���T:+�\�?^�Ξ� �8�2Y�$�<����+���X�n�݌���d�˙qIq1��(���M'���F1�K�������k�z�'}mo��<l�3�vf�N��17��q���:펷97QY���t ���{V�}���<��2�����lΤ��-�&��1����WjT֪��FOw/��2�!�,��g�!���7���x��e���v�!(.뇱�N���4Zd��c
����궣;��ۋ�ŦM��h�>���*�Y�in��.l!m.��������a�-���e.���eD��1c��w�$���;��;$`�E��#;\*��&N����0�wc�fds�6 �R=3�6N:�x���G�y�0u�����u&�D�hwۭ@SS+n���ev�O�D���S���7ޖ�~�Ǌ�ܹ�/���ǟ�5|�m����I֖ -C��� ��y�bG�5*i�����u��Z��"�?_�-�*1ϥad�(7��+?\�-7`���	`�n���?*�ɺ������w^C��=R=�κs�3��9c�����.dhl��#7r.�$tГ��Ї���?t��?����}{�����}@�7���Wm�~d�sZR��B��$�T/��ψ���톟մ[��Ϊ.�ģ���G#ʜ�^��o�!������q�89?��4�U� Nt(Q�?q�-G��1ӷLi!��(�EE2r���1q�x�5�S�YVM4u'Òv�$:�׆Tu"�A�LNZ����v����_���<���e,��t�·Lq�A������g4���Tچ_�	�-��W�����?�@�A/�o����{u�"Jf@�����/����0j��w�xq�����1w�<���꣩�A6��zz�PR\��#�]<ދ���&�^&<˗)Q�Rq�3���{���>Ip�����d,��᝹���s�e�����g���\O剠�4|7f�M�;E���N��������{��ӧհ����x�w���U����,Q��]��-<�ģ"JD�DiIN=�4�&��K��'#���Y J<�LH۟:�ւ��\�6>Z��`���K.�(����mR�{�	Z<R��:����P����$z{�;��n�GM�SϾ*:���n8��J�)�6�e�V�:�v4�j��!'��\��q�qG�G̙g��:$2'Vk��e�>ukp�/~.	�_�|֭['���t?�@|�|�$���/{�1���Kr��1k���u'֭۠F6>5a���V�G��JPO8�h�蘣�r�����s\A�Ao-~��[*�
]t��ܸ��kQSQ���/C��ZlX��E�Ǣ2`'���\�,B�h:�^C��Q؛�����p�X��"
&tbjĽ��x�b$L �ya\�Q�5Xܿ�΃����.���s��m���>���oy쳆~����-���ܤ�tR�y��C*���.kn�R`����]	�GG��<V�ܗ����âP7�2e�.U�T�jsv�@��n�j�(j�3��fB]Z`�1cp���bP�����S�R��8��Ǌ|&;�B�mIC�J���,�xu�մYN��?���q7R��3I(�!g@�1{����s�M� O�X�|�00�ꕈl���I/�}M��gh�A�M�_GCsf�yV�%����)=�/�1�����/0d@��'��H�H.07�-[����x�di�lH����^~�%twӴ�������U����:���C`��ȫV��.w�Н���;�|��۩��R�z˝AO�gqi��<�K˔k�=�a�D�����Cgg�h�s-]r�%(/)� H4���ťX�n=��aa00!8��q޹�H�����g�Ą}ơ~{�UW�왂,����uR3EH��	b0��e D�������+d�4i�$\{�5����7��glڱ9i�H�����{��3�j�Ǹ����%�H{��{�Iº���lI�؅�-������o[Gn����;d�cM=ng�|"~yṘu�C�۱cƍU3i[�W<�=.l۶�D/n��F�ji¬;�B��FaI�y�8������oH�}�QGI@e�kr����w	��������6��{}~��Fo�ޤ�:G7�&����a�+W|��vI���v'�7~"��7�^��^z	�[�؅�?��:�9.}�7���W�(�u^�O����l�Cv�A#�c����8�\����{^�pmcǆ#.��g��-Bܰ�k���=�l�{9L�U�L���]��7��-����W����o\$'�?�����i�gS�%�`d��r��� �%��l.)H��H�vN9�GH�2xf�<���"l�+[]	�+��:[�l
m�lV��Ga�@�7L�������d���X�Dv���]6�,����B���fTx��,��bW���l���+W��K��&��:zz��%x���ȡCe�PU^���{�(+�t}��:9t�M�$� � ��*`�aĜ��3:�8FF�QF�9�QI""9HΝ�9}r�o�wW�}�ݻV�{��8ki�O�ڵ����7N�ET��烬����NfR���&%%�A��t#g���	�W˭;�����a�ƍ�&�9ɓ$�\*�i'M��o�	��F�؂:���X�����M����
�}yH�sp:TB���*�WG[�l�?|�������LU���j�[����'-o�M���ժЕ
��WZ���,�Z�V@��@����R\vɥ1|8� ��	��:���v� �@�y �����'`HV��^7U�$|��1�b�O��~���Z{�w���a�a��~������Ȉ�뇝"� <��\nV��q��-�n���n�)#���G����ʪ~�ki�]��{����S�JR�C��N�������p86�馿��3Nƛo�'{\��T��g�����9sB�(�e�>�`� ���@�ǇsN���^{!�9�	�_�@�Wԡ�v�Ka8�i_Jz��/���۷��9����Qf��_}-�_r^}�u	�_|>^}�-���k�䰻5���$��z��2���NЫn{S��}sS�%��o�=7\u���>��}��4#�	n!��c���������ԌY�f���Q�p���=�|��W�i�ؾm�

��wt�.��x��FY�k]Y�Vaz�x��uX���o|߼�e��d��G�X�)j�6�G04����U����1#G��ʽ���[����p��>�$���֊�?����P�DjM�(b]�0R1qH�hv��Rb5J�j�(���	&��3ϖ��o���/F���a�����S�����i���<�4+�ʥ2҆s�2"(�j�@�������,�1��o��9��2si�ї�/I�p�&x��ie_+�h6'[�:g�-�2e�P�ަ-�~�n��y��M�x����h����&���^�H�._h9]@}��p�r�pb�������QX���}�����X��gq��&R(��#G���l�E���s�X�K�Ȉ�g"bw8%�Q&��9����j9�.K$���b%��#���4)k�B&lJ�]�ڤM�z�*t>�U}[ �Fd�J���+!��,s^wk��Z������wÆ�K/����::��� �nw"�	8#P��fv&�j��Ȫg{:M���C(�uG%�o.B"��c��믑�1��/���9t8Z�3
J@g=��c%����- �±8��B������w�n���ŕ�\����`�]x�����@���e��v����*�J����	�S�����ko}���v �RA�`���p�o.��t�C����N�[%�{}����q�9���s��w�)�:戙�h�s�Ϥ�R�5�x�	�s��y���&�{=�~�E�=x饗d]�s@p����W�]zŕ�
v��އ��V5^�#C:�dn�t#��K.ƹ���7^~_�%b�̡(D�qAM�@�~�]�'�r�77��C"��7���=���0::�dF����ڮ$�ͮ���֔�J�֠5O���ޠM1k����c�(O'%��D�Б��!�����f��ڡi�_Y�>��7�t߭�q�X����އ��C�k�=���onk�>)���̥�u!	 	�A	U�.68�$@˦I�΀~�E�!��_ķK� ��Q1� HLe��V*�t��fec�윳:��\6��g�N�U2&�-�O9C>}��叿�N�xL��Y8�&m�._��Uѩ֩s� E��H)��E�bk_Lgrtq6������%�����A(���#��h�[Q�R�|��2�8���E�*n��N+]��Lo(�I0���v��_?̘q��K����|���z5lT������8�Q�s�i�v�DDm��M)WV�|�<��H��B����~5��{�n��lomV�f��̙#��|pӲDW�� �B�������W���	Z����cal��zXr�VKު��6��'S�����	H���KQ�ϗvi{[�s���}�����$�ae{�Q�1@��[ I����m�����D3�K*�,@�m[7#����|Q�0$́ѣG�.ej�3����عGf�L�t�����;w��p!Opo��!ؽ��X�Nc�I�te��dA�yg����:S0"�se dg �H�g�L�e�/^}*��':���W���ǞDw<�h*"��9�gL;g�y^~�̛���;�%��(�b2?�����/Di�_p	�1���������^�ܗ    IDATw��E|��^v�l�ܭ;��F8\l\�[I��0z�G;�p������.���_��O>@S]=\B�����O8�\{=�����Y��9:��|3�L��7_}M�����w&���Jjb=���wﱑ����[�P+r�n�*��)l�x��Ƃݍ�]�М��B:M��U71|�5/����}܂�և3�?���$���F�����7�R��H2�x����n8�64Qk��X�:�����N�{��8�䓥��ڻ��ӯ���� !��j��Jι1�Թ��U#��V+�������XRi��؍\��S���[��[sE�홧��g�}/-��&%���!FJ��# 3V�v��gx�����8��Y�0H*٦�i�f2
�Š��$x���6%�o���9�o:�$p�W�����e�N(\ �Tl�>7��Æ�{�EEu��B���X�i3bi�R��αC*ڍ��b{�h����Kgp�kSP%�6t4.���U+EO&M��ÇJ���'IE�J~�����e=R��w�L���s�Q�5s�Z��1�l���;�^LE9K�j_Z%ׂ��V��ԥm�R���퇚�*%�cr�[�ڤz&қ�g���ɠ���|�>�ʫQ;p��`�]� _|��$mtO�r?����[��!#�K��N`�^�� |~/�x�i΃�T^A��؍}�2?�+*Aye6o��V&'cv�HC�\ęU�l��?�T��()��Iq�2�k�ZwoC=��f���8�L�py^�<7�[���[�Z�� �ҕ"K��񣼤cǎúuk�/�� &�"֓T�.��I�L�Q���C�����������Ԅe�W(9Z]�nи1cQV^"k�C�e4���6c��hm��_(�X��5�B�h&-|�Q�?\-J|�y�Z4�C~a>��A����GK2������g_���Q�Zo��fL;�|���hkj��=��������(L
���HQ笊�R��(����Q�I��N�w,V���@)e�i�	
�Y���?I����?�����������?�g`@��I�
�>���O>{�%�8.��!�B2Ў\��t
*#1���ȕR��G�q�)���9C��w��������n��g"�%*s�&��e;�;���,4��ۖÙS���?�=QW���CX�lT��6{<.矬��N���%��׉<�D*�I��%Z�7uUu�
�n��e�)*,�p,*�jͮ!���tР���H	z:%N^��$h{ҩ�XF&�QL�/�Q7%��r��6���f��_1v�u�Ė��щv�z:���P�x��U``�jI*Xe�R�y'�*�NK��ܘ���u؁��Z,Ɗ+��:t�T�˖��_60V�ܔ<�{X�_���
�<WJ�L�Yhvv`�-�j�[`H+�[�$|&(΢1��1 �w9"�	p�����wP�]�����0
�.D���?_,>�A4��K��׊��|oR���'M9���@"�����nI���Я��4�!ۅ�0+�n�S굠����EML �2��x&+�E��rB�!sI�N�i2�f"QNԾ�K����!��'�6:ߓ�������3��|�'��D*g�c!MXb�,ƍ��;w"�(�$�2�$v�� ;n���tJD�<�"-o��8EJ[�e���T�K�k�3O;�i
Iq�fI��2�b@����~�p�{�)(��"g���Z�vZ���f��x��O��܊d<&�0�w�q;�;o����E��=�ţ�]�ho�sf�G��p���N�;#����8KJġ�{�Lx�Z��ǁ��P4{�R�n?2�0;>"a��0���cƎ�Ã����>n�������p�xȫ��~O}��;�iǱč���jE���T^
w(%3�,R�\6E~���.8�t�'���'x�ӏ�Ѹ����
��o�j�~(s3�S#����$���J$2���5�$��O�K@�x�'��O?	�����="V�V"+՚�C0���d�ݸa�CQ����Z,���¤4u�<��@w h���Ê����-�A�
��`��ަ�_C�2��������G�?� ����Pڸu�����ܢz���ѯ����b�#���-�DҕA�M�����KH )?܄���6u>�S�4���ԑN%�UJIJnfl�9�@�b�2�7�5�Vx�޶iq����/���g�b�@n�ݺֽg㿮Э�n��U���xT�C�6�Pt/�8b�̕��RU34;��Mq�afɊM4��!+z����f2I[N���NtG�@�:�,�K�f����W_�CSK⩬T�eU5�8D�j�Ȥ���;���0���	F#�����<$"1�qM�<�ƍE���$��Փ$�|�����H�	[��BaA����kk%P�"W�i'M��C��4�i'Al�dR����N�J���~b�jΔy�`�G\� b�4�a�ݼ����X2��FD������Q-[:�B���K��¹3�p0f�A�!
c�}��s��E�����pҤIx�7�v�J�~�C
�y�۷��7����@Z@8����FT�ĝ�x>�5 BW6���QAm�LB�n
�
�:��9�HR�\t�@d�৺�l��F�4b��Uӎ>Z!��?��g`@��)|�-R�ܻ_�Ӕ�&��@&F��F�](ln/
��ͤ����HF���$ߏ)��N?�P�}�	>��d���ܼ��m�7XWČ�Vl7]HU`�a����f@Ϥ���q�d��׊v<iO<�$���{��JJ�1��cQU^��&~ieJ**Ek}߾:�Z�^8���Co�h�?� \u���YQ�����f�l��<�b���5H�U���|��[� ��%e���?�}��E��C&�C����_{�� a��q��w������1�_������3�����G� ��;�;���Tr����2�(CU�!͆<�8��>��C\�d��dDΒ�}_Kc�e*������y�5_ע���������=k������&�x>��U�[��`�4�)9��}(��&U��crE���(G�T\i��Š�'�.��&e~��F�{d%d�T�k���d���E�9&KT9���k0o�<��Q��|	��Sx�Ï�p���磰��ͭB�d�EcBe@����H����m!�k��`���P�G9w��.T�� ϫ#L����Ģ�PSL	�Y��gO�9�J�����U��	eO���L��J68��g������$}l�1$��!Q��KM�ޟ	&����cq�\� �?�[�`P݆(a~ފG}�w�F��A(J�x�C��;�x]���iǤ�A�~���A�啀݁�6lĻ�/](��3���kp�y��g��O?,��|��{w�@,��(-��Չ���Ny���S���Q�p�Ǌ^����W�����c���A�&dv�ਸ਼gw�Ќ8NHg�^�9&�ኲ��tO뺳d���9��]K�Ό�ш^�ٲ�l֦�l�]��z&����0���r�\ΰ�9]��9�-'?��6[JӴ���i{ƞ�:2�\�e���rV�e�%����dr��s����TLfs�����z�4l6���Q٥��� �p�\�0����%���i��%m)ݞqس��۳�lְk��g�
��k�tFG�T�t�x���\l@�c@�(*������ٓ��6mM�"]��R�Q<�Uo2!#*�_y.��ܧ�u�;�x��w��Ws�aF͠�Vh�� ���_~im��/�g�j(�{.����&���]'nL4>yꩧ��A���]x.

<�,-BYy9
Jʩ�&sm"`7�ۈ������E��?�lZI�z]��C*��rV->��MO���D�.��b��|��ױr�j�V����vN�:��>l�y��>g�L��m��+��ȑ#q�]w����a̘��/Z"�9)�hoJ$6�Y�3�L&ϏjG��S�k��쬔��7~���f��a�6)x��c�J��U�+�n�&mʹ�d��k��um���{F��{	�浴��_5=lJ��:�[Ǒ) `;���O>��y���W,�.U�˴�̤T��5�X������*�:�	\���Rb�$##�Vs��z��)H��8�_e�����6|��W�9=��WX�}4`�x�b�RZ2���!��-M�2�9))��@+�#�8��v�  ƌI_t���5� �Jl�Sj���G�5����+V��ھ�Iz�c�f�B���'OÌ��$��<�\*i7�i6��=+;]�"��T�Jƈm�����ȈϺ//Ox�-��9�,^���N*Y:*x�69�6-�������	��y�,-\��4��/œ�>-��<?�X_t���<�ԓX�r������
J��h4,]~^�<���A"��Nr�P����S�L��i����:��@���H��$p��vg�Ԅ?�~`RD�����9;�"
ih����!��1���h 2@�*�L��fP��[��в��4�z��\�٧DT״��г�8���f��0%<�
���iԏֵ�-��Nt-�BES��$σf�6C���c�t]K�9�d��C֡i����	����s�d*�kZR��v�cQIa٧�ƌ��ǰ���?����}0
�|��k{��ӭ�jn�	�o��~�]A�RY1� ��E��%�2�v*�ۂx󭷱h�2�Hcu���+@S�[=ԥ���T8��!:r�� W6	���i����h�x/<�<�Ν+weE)���2�\T[���R�&Xͦ����ѡx�۷�D$Ƨ_|�ŋ�P�X�ћ�� R�������Ya3(��;m�4\v�U��������E�ɚ�)�����������߰��?%��}7x�³-�(A]s �?0?,_	����ō���%kM�y"��B�����јTՌz���|�n��MG$���'���W0G�ԅ�L� 9�YЭ��%
c!�-nz�klm�V%ϟ�v<��F��
���.��h�)���zl�s����3]'g�l��F�gV����2 ٮX��7�֨��M����%��!�D���"�]%4��_#�Q�	� �X��Ob���d������E�]�T=5b�8����^����6��~��h�~�H�w�?p�%$ �n_��޹�8�U,9s�jy��p�,Z��6l܄���@���3(��M��c��
�r�T;h���9S��E�c�I�&�X38c7#�	^Α݆@G+J
��!�;�C �̇ł���Y�����"����p�x�vӟP��G��[�垝{D!�H�[T��� 6o�!�~v�hfs�y�J����a���"�D��t:�[E鏟Q��l
'a�I�#p��E��3���U���LDq�q���֌֦FD:;��!�dm�	�8� ��A=)�p�I�eg+c�r׽�bSdʲ����_��?����3��fo������}�馕l[	��vz����]o&@ﱛ��L`l��`�k�9c�nl��pn���7s�qǿ��5��������`�u��)��"�j��-�W7D[:�4U�Xyg��$��~�8b�(�_�d)�[[��g�J�۔�t��nv��c-h�$gJ2r6�Ѥ�p)I,�8�X�t�U�e�x$��^xI�ۣ���_s9�W���_� ��l�r����k�BWF������{X�z����R�,:���]]]_�{�����yy�w圝���?ߌ�G�Ǧ-��t�
#Q���;:QQ���U���E�y=�qr��|�)Q�br<x�����QTR���v�s�X�a�ۚ�ƤY3�{5�]<�ܬ��*I<�e�����.;�dr� �$������c�#�a�U�u��=DX�J&]��p>,�XS�j���SZ7�5���w��Y�%�������pX}������	�b��t��8�9M9(=ʀ/� 
�������H!g��0�Q�>�,��� �w7�҂b_�D�-\*�)��.��X۷nC��C����'c�����oVg��2i�s�M��r`�A��+��@X��)R��cp%4��v�5WȽD�;�阋�_.(sv`x��#8�X&�4Xa�O���dR����!x���ڵR~�U:1b3*��r;�#��z�Lj�����%��"%�M�����cp�o��tES�9{��fhOO,ߧtG�uAUeŘ���{�H,[�XDl�M9	˖.ſf=,�IIbQ�2'�����mǕ�_�I��ￋ�?��:+�E��{�v����e�Y�\���6�80@�<'LD��`��Z�V���A�L���z;�ˡdbr�����w	qlC���&4Zi)
�RdϴQ0+��̶�u� ��}�kԺ�z��,��_����ֱ==t��Za�±�:���a�;u�y����{�;�$��#�&�_�z�������#�;�U�/�zO�[�P�3���!bL��p A��=p��0�x�N��-`v�تd�0	ɠy��4����"�!�L�؟ʂ`�05��=�3;��d���^�`���*��w gM>7�p���X���=.��2\}��8x�A�ׯJ*ZjMS��-'-S���\�RZ{Ͽ�v��-3�c�9F��wl�%����DW�E%Ţ�EyɃ���\�)�N���{�n�z��uH�!�����P^�W<{r��^�=yx��װj�Z���eϞ�(���b�z׽3�f���������*��y��+7Ij�Q��M,CI�����/�ǥ�9(	(b��"6����'
7x��KT+_9�H2�k�kɒ����Zv�2��_+o�w�:ۘ|X(w�
��0XZ 3'q13g��k���1�nW����<^���َ�mBCc@g���!\��\B0����-)*��(���:
�]}� �_}��Z���b�+4�HX��]:�tu�#����~�N9��K��oA1<y(� :�f<y��⚫qԄ	X��R|�����T˝]�HX�RN�t���Z�a�W_���ު5��&��9
��0[�V�����0-uUg���1T��k�)3޳D�_�k��ߊ��5�O�E���/u��(G����Dzv�K&"8e�<���;k�J�'������$C�=��y��3O`pM?|��X�f-�rӟ��o��=�|:
]dV��@D>�~n��ZL<�h,��|�p�r_�{Q��a����6�۸�����FP��J ������{�,4���0t�5�q�t�4�"�#-|�gv���t����$i:G��ϿM=��AEI)X���-��*l���`�_�r5v��tɮQ�t�T]=&��7��b����7�)��bs���l�S��:t~T�����yg�2�L�;���5�6�s�k�����^Q]}���S�0�}�N��?�����|���6Ƶ�3��cq���hk&�vd^��)F��cT�eyR�TA�֯݁TNe���%�X	>���̗�y�tTU��3EEri:����3��υ���@��X�`Q�P]���C���R$�	�u�*X����UӰy�V�|^~�e��	n�8y��<xȁ��ƿf�JQ�z�w�9v�XέJ��'L���{�b����DB���JG6��|�D	���;S��e>��K,\���n(�f�e�hl��=3fb����<>iw��ޥgz.�Q#�������*U�wu����w�??_6���&y����f��MY�pQ�����Gv�P�֬Z�6��6I �w�����fUnbB{2�2����m�w- �U�+�B���a�E�
�|]>�.��7SY.�֯�&A-���͓J�:��o�������z ZVdn9v�̴3�-	B,ǹ瞃���[Ip�~�9�x�eQ�	PUe)��ރt"-�ᡇ���ɺ 7�t'J�nڲK~X�X�@Ye��*v��'�m���[o�Y��m;0{�ر�Ni�s��,*q��k���-���v�"˖��CP�*X�<���b5h`��K��� ��h�����Y9�L��nJ֚�k���,���t*�uQN�ipI��J7��q�E��t���f?(yF]k ��d�    IDAT3f?�%+�
 ������� O��<�\wťH'bز�g�}86l؀O?��P��J����&c&@�x�\y��,}��X�b%���++*�N���=^Q�S������%-wޟmmm1b�0
�3V�l�1�܈z��E��M{�J�N�'�Q��x?�� ��P�;0�$S��ѩ�mz.����#��A�leS��3o�!�#����]�#cph�KP7�fI���us9ͺ'���Nl�7d�p���?}e��.�<�+��r�P��	��emRV���ܙ��|^���[ϓ�i:�*�` CoMg�Kkzv���~�cX����x�^o�V=?�ۏ�����D�5�CtI�er+�df'�\���\M.e�-��T�\qĳ��"J���]��/@9ڍ���c��,�$�Kv�8�l���4��6W_x6�$�����cذa#�\���o�(�cVd|n����# (�jnݼEf�/��n8�O�,��r��G��u�q���KYaI1�x���Z���^+��\�v�K�j�+e��K2�F��r6/��_�V������!Cp�]����M���l�۶9�G�[n����M:Ə���U�)H����u�蓏)�'7R[S�TC6͆kQUU!���83$Շ���a�Ŧv�ҥ�A�͛�r�͹��b�-KHct�-��y��ښ�j����A��ằ�pֱ�F67U��lV��|mq������KY\V)�G�8�����㥥Z]U�@[#B��T���,�[���'���믿^ѹ_~��^~�~�^�U�����mR�r����!�BEE� ��.��	�Y��x=l~޲���p���w��"�{�w�}*��P@<���TWV���[v6�;�A{s�:e2i�	��T�r/�mZΤu0� R�Dm����B�	8�0�/9�}nUsL�-��� ���3�%+<I�Hus��(�nc��/���\
�:O?����κ&<��X�i����V� 3�t9Ԑ�qRx �M9'�0���(/+z�hI�h�mO#���C�;e���?봓q����>Ǫe?J�N�&�I�67���	Y�ѧ\}���&����)?/�R8G~�܋�7�k�qa���@;�ZZ囹�3�^u��R��2�*�r�R�g��rݮ-t8]]Hg�4ʵ���岆�n�@�f��a�C#Z�l��˦���5Ùc�Ěb��{Z��5Ct-�Y��tM�횦��ɽ� t� 1��=����D7��r��Գ|sPO�	�#4-��z��q���q�5�Me���ܱU�&џ�_vW0�6Z�����'���;?����x����$�����}|.d�Q�c�ht��)�����I�*�~ȩ���oW8ge�$l�����T�T�SIm�=s�^:�-]�Xq���6��~�4\?�83@W{yx�l�&<ރ����C���Nj7=mI�#��Еd�mع{7�{��5��,�.R6n��͛q�y�a���B�c����QQY����˹seFw�����K@_�n���4Xfu4Q!�U%]w#������aņ�{�4h����Jʱw_=y�	l��G�N;F>��<��cHr6�N ��'[��#�(��?iz�f,����"�L��XcX��r�X���q�H�Z����`P�i{����Z�V@��jֆ�k�Moښ��̠��3�[s���7��� 'N��*�h^��tF��Xm����i��=�yO<�Dyn��4��^���C$ǜ'��v
�$�r�86�k��z.^x�YyVQe�hmiB,��C`%`y,[����;�Ņ�d�N�nF�<������x@�D0�o�+v׷H�v���/�?��+�C!�]~|>wf�y
��m()*��Ï@S{���٪��n��SIL�x*�K��H�%��L��f���x�*���{*Q*�� ��}g�?.�I8�Iz)�="�sJ����� 6����Ç㹧�|���f�|�E�ظ��� ���#
��t(���� c?$�3ð�������;v��_
�=�"�����﮻�>��-�έ�JK$k��'�{Z��'@7SĊ])�K�בk�םA��#?��z"�"!��tBX&"��Ӎ��D���C�yx�e�I�����|j���s�
:sl��dK+N��.�3�����%��wk�:��^X��'���'�{�y��3)��d�lְ����ެ�I�r�Lư�e(�բ����1��c�=����������}��g�5>�u�u\�(�D:��)d��>�A�C��0cd2�����8�����K����x�^�F�^�d��i�Q)͍$U���`tu��j[x���qӥ,��
��
��9� 7Tr^	1bZ�&�8%�*�]́��\�i+j���r�?t�Kc��S��K΀���s�<��˗��v ��~>�WW���Bܛ�JlZ�[���ۺ���Ė����R��}��G27=��DY�k�c
A���_]n��o���<�6mªU�d�8h�'c�FF� aP҃`,�>�?���ˉ��o�*+��{�>����k@��Z��H"�����A��v���i�s�I��R�W����@gwX:���u�V����;Ď����oK�.�m�f���hU��5�����LƬ �{��,�D[�Z�yi�ӵ,U�;��
������Ce\�cw&L�����ض�ضm۾c۶�I:�m۶m��=g�g���jͫj͹�QQM+�����M���X�%9���{��?�c�v��#Da�ɻZ��v����i��y#�7=��=B����Κ�׃8X�`���}!���mʿ�GG%�F�Z{�y2�v�m�(�@2)��gq����7]'rЗSUt�_/��X��O�5�Oi��e���{uyC��Y�!>���s�'Ɵ�#E4h(������b���*�����R�2G�dӤ\���i��r!�߀��*`�J�q�t���^`����*MM929H�u�J��>����v��+؅�6)��k���s�������2���#�w���[��|�ܯ.ܛb#�xW������Mr3��ցX�T����y������U�ݤ����?���+U��`�OO��풗�c����r6:z�����#C� gH�pI��",��`�-�i١�7�-�\���bv�G�L$�<�ߋ���X�߆�_a_q��)d?�+� P�{��)��S]Ԇ�h/;T�kU�Tt�����l!k��օU5	{��Vʳ�K��)�}[m�v�
��Phr>E����1vZ6���[6hN�ǥ�Y�P�����?�=�DC%�dyt�-K봌�Z񰳲n�J�$E�ai:�6��d��¢q��B����]�.������7V��>����pL��ˍ>	[�#���(�q��e�u������ym{�8 Aa�����B�^WD^.ȍl$c��ƾ"s�C�]{�OPo��#�/pe�ik~[L��H��I�A��%�{�)A���E� "��Ll��U�����Gr:�8� +p+�w�Q��%�m5��^��.���҇yXx���6G�8}VC��*�^�0����]��L���k���,R�ب]IK��/{�jv���藄&�6nLx'�Y�<В�J��kyin�EM�bb�}wnE���z���骚R6C� h(��Ϲ�����aP���Ա�;klN����IAM��!�|�͗}�v��W���vDǍ߯�e�D��K��u��Mu;X�n�7"�usc�P��"&��jQ8KmG?��)�X]�ĵ�鐨
��6I&�LhD��JT��}�C���?H-�ވ�:�����n���%k�n�M\ॆ`5����s�B�V{��Z����K]i�d0�=CR��Ӏ��l|�:s0!:���s����N�Jȣf�d��a��v����Ք:��K�g]yj��6�@��E��0�B�럣���}�a:���?3�/�ܔZ9�䢃R��UV˅�{��c��t����-K$�?u��S�X>N���c�1\P�Vl��܃�yx�k��>@�������B���\G�x�_�巑�)��+.t�>m��稊���'�Z/��r+��q���l>M�op)(�B�>锁�̫�H�P��F����w�v�Y@)fs6��{5tқ +j=�h��|Ey��[��LDR0s�H�u+�N ��݊L� |Ʊ� ���M�긽�Ş"����v���o���]�c�a ^)��`�,�aw�+HI��>[��C�Fd���3������Q^Z[�-�kHz��m'�h���ʺ;7���*V�g�}2�2����b����%���C-�i�+B�X�J��	䛻����U�����z�4��l�x�θ�v��Q�Hԓ'Ci)a�\p�_1�Ѐ��n兹*3z�����.`�R�����o$��P���. �M�d�w�5R���I�q�~���Ǿ�>@����*!�O���]+-7���}��eGTX9�rX���Y�}�5���ʛ�csat����`p6��� Ps��/o�ؔ.��R����p��-$! ��~�-w�(f`v��s���"=fXώA�g+�[*=� ��vy���a���L*Q@������� ��wX�%�- h�v�I�w~TҘl���1��$��w�t��/�0����UR��2F�<5W8]��ct�FF|��L��o#*й�{hB����#��kvX�h�x�a�ԛ>eg���"q��mr��~��,��.��߅�Mb�Ń%�Lk�{�>���DUY��c�v##p���T��@s��M�Z��A�-�j�x�� �*}�|��s��6�;�~Eu�@��D���@���c%'��En7�y0���v�Q�N���Nq���4=U%�Z��[П�q������T�n�[�Q�g����elxyi>�ŋ[��c�F�T���Qbfh@�8Z��o^�>{a9*��>:��(cx��3�Y��+�h�I�?�U��j���dK6	K3Wv��<7К��YF�q����j�$9���i��<l�%"�B�X�����Ԕ,PC�+��Nx}ږ�Nb�פֱּu���%7�8��o��O+��j`?O��7��a���g/�`�ND�������-9����78�%-5�C��T�L���A~B��_h0��ڪ���"�����I���ҩ�a�u�(]��f+�߁��h�B��X��(_#`DJ*�����av-����	�m+���9� �]>�>|>eɷ��L��{�{UK0#��'����Nu=~���&�KT�V��X @�%��r�`O�Q1�һ����ϴ�#��%|�ʼ������	l���[����Z�7��VסOtީfm?���E~���9D�.�b��M[U�j%�ŵ�_+M�Sͽ}n���6a���0m�WпL�ͧm-�@��ޜ��8S�e�����O�i�#����[�IO�L������V��EԄ��:�b[[;Aq��Q��������_no��ûҪ$�v��Ai���q�(u�K�"!Z�ø"���[\�O,ϳX��Ⱦ����w��A�F��4�~��"���h{�p�r��s�u��)��B�F��q&5Y�T���Z�!LzI�<�DjN�x�-K�3�W�kQ� ����h���=	vXI3
J���M�fh�"V�jj�S6��$Z/�k&e���Z�Q��^;��<�X:��]L0t`<q���tm��b�m�_��OϏ -�����N	x�6<��(��EKr~/`Z؊r����5g�q�����u�����k�~ڒjE>��	Ov��4Z�$�µy��J"ɶ"R�^���ſ^��o:;NV.��4��U���l傒$�F��>͆Q�䓑�L+�i��\[;K�|n���I�zM�n)N���f�5ҫs�<5�ҮQ,0�!��S*	,)QT;�!r��3��9q���3cDw�[C�1b}]��%����R�Q�E�-g�_zel�Z0��p �=��^�Ў1
�47�m��|������?�A KX���jx�9�)#��B -(5�=P��4A]]E�i��1��80�aq���f���"�TvL����%;1�lz�֚���f�.�(ZS���ĩչ���kg]mrD+�R9����%R�� V�Y�Y� ��X�ݻ���	@�^EE���Nsgc�S��E�����]j�^�n0[?5�+	R�@(�h'�������d��E���V1�����n��&���k�ɥ/E��E��s��[6q��2ۤǭ�j�m���s�7�I�SbzJ������b�����~��4�W��0}�5�G_�	3��iSָE]ٙ:���=<���C&l�"�m�	�JZ��t�]�L���z�vp��mi�7��P�>��3:y���j�;����w'�^�В�#���Í���91��n���sMOP1U�Z�(**��,��������@%��J=lb�_�*G󸳗�^2"�$^���;�r�F��6;	ڥPv�o:����:�5,哼c�G�6���D����tS�p��|�l �3�S)����59D';�D��Px�8yK�U������������g&����� ���w�N��[��;�+=]�-x.��@;�%������/lY�`����������?*Y�����͘��fga�ϯ,�@�r|{'��S�l��	UgV>(Z���H�/�j�R�{0ɩl��µ̟�t<�A��(�d;sT���ŕ��}��c�KW�S�c�C���F��
J�5�'q��=���-f3F!V4��$��C�.Bێ�ϤR�p��Ǘ���Q� �_�>�w#����}ӷ�UR�i�c&C�َ7|�xO�Q-���
H�ʨ䘜�F�bP(��k��L�����T�/AK?�d��))]d���1B����U�$u�Hm�P��`��t��u�f�//n�|���z:����V���!��Z��W�
h�	��?��\y�HNĜ��-�P�T��g�8�&�������(TnC�>��$P���R��81ʏ���m��n7�C�L�j��΄�I�O�_lZP�8���M������a؀�B��>�N`�v��	އ��"Y�4����u"L{M0�uF�; �c�\��n�2	2�AP���M7��lOrO��o��J�V	�P6���@V-�2�p��@J*���4��g�)���Z�y'
Q�ھ���h�yN�ϗ�[|
ˈ4�`B���b�Ki#՚�pD��j�5:�vDS�;��C>7���"���D�U�d�������&�}�.�K���40�	�_ʌ� 3,T]-Q~�j$y��v@FL�;U,���Rti�@ F�/���x�}J����CM�
KE�ld��qߡ	)��)˜����ge!�xm^	�5�̳60/��UY'2�]e0�-���vH���`P4�'�~���@�@:wA|�xY��c��`n���o�h�|t�H�#WB�K�mx�*j(5����v�:����nЀk��n���G�p6V{�@GR��	��Ԯ*���[����w�1[?���%g�4]��
�8!�i����z�I��F�|�nn��
�·����zu�K6�P��_��uk��7@W�TË�_dپ��8�`�X�'s�ijO ��2`8O��$�/'m�hݷ��wtC	���E�����_/���S�/{u�#�tHӂ6X�t3���pM�O:R� ���SXq!���>c�Ԧ�P���*i1G�%=,0��r�q��DĆRuh5F4ms۝N�҃^�X�fnф|���7�����j�����b�ҡ�[�,>�Ӣ�y����)5�p	�Qq2�rC9���L��~���p��ys��4?�E��K�`�xQ`7*A	"9u�V��d��#�D献��s{mi	j�_�/������'c[:��/w�4����5�ۃ�#����c�]*�K�R���˾���#�����zw��`�@ɇ���%���4t�����I�LZ�P�r��8Q<���Kg��L�'c��ET!�1��U�s���N|/��mul�Ȕ�&OEN��ة�޲�}�ad]�;���-�Ϝ��o;�t����x���S�o��`�rQZ�8�Ab�� ���Lv"Mأ(m�B�Q"�t�n�?�N&�e�{�z�	�o��=�����n�nLm
���g�K�%+�%N=��ߙ"]�F�l��:+�aV\�v�T��
:�F�|Ԫ툯oK�� ���K(Nc���5�k�<����!h��
{ڃ�D<���9L10����,���Gu?.�͜��ȍ�B�W���E��_$=�`Ρ��_V���:.TP��P�8�&vk�}����W���RMQT���G�RI�1݈�X�(�0���S���ݯ��X�m������L��q�H�3�N�7*0��%��n��Qr3k�����qÑ8nw�����D۝bwJ�x�h�#j� �5�D���O�����	��@������р�s�h0)��R[T��?ߺ�>�\1z?�� C��ٍ��"y���+�s��XR�(�ҲmK.��)dֲ9�x�r1#z����<�u0G�m��|�`�?-��r���?�ֺ��;�J���2���2��Ño���9&�!�2�?ݞ�t��Ziܦ~�,�Ԃ��rjT��Y4W���)E��d�Ur�.��������j�2�.��I���*��{�ހ�W���Ŏ�NC��j�</� !̬_�iuDD�f�;����Ϧ������w⑀I.1���j'0��uR�sb�^(��?\�|�)�}،�}�A�~A���jbʯ�<�U�����)�k�dF��{��+n%��z��h�4�N�P���B�?h�@�'{NߐH)46��0���9"����ĭ]QS3���[�
���D�UWL��V��fp�ꥐ�OM�y˙�2]��=ӭ���Ft2��O4��u6����b�2U��p�Dy2ieA��Vz!O��	}J>1�D�A^�ٖ*#$)K���.Y�X��(S���4��%����1���dm����zT���ـ[(Y�֡�'ʫ��;�f�ㄝQ�N�6�EL��?���e�՘�8 t\�i��w�
�����k����"������'���Us[����{!!���W��z����D/��r�u3�ܳ�fd���/2�U�⭷Ս���P��_� �?�E���h�
(���t� �X�T�:���A�[<�i������9���e�f�"vTհE-�G�
&V�g���J�*��TnPv&hrN{]�����T5˷G�������4�r��*Iq]����h�
�������ȫ%D��@��|��nz� 'w�p��S�S��y�b2�s�b+���x�7���Bm� 6ɅC��!BM�y�v`@H� 0��4g*�N߲�

���T��s�q���R��O_%���X�u��w f�YoE�����RY�~d�cn")�I5��.բ��iU>�T=�d:�N�k��%��aW"ܔԽ8+����v����QÀ�M��U_HR��0����5*1�3�c.]��.����Ȩ����  q+T�Z\Y�A��	��.�Jc���9١׍]��*,�E�wA�o}@8c�K���	q�v���c�k���儾���t���:��D���>k=m,���W�$E��_�@���S&vS���o��V,�`,�h$���"CJ2D� /FS��= ���9IE������h&�ע�	�H%c0�}�+QR�0���g$r�9H��=o�Eu'����P��ۦ��iTۼ���9���F�K��(�B�ѻ$��hRC'l+_yˌ�)�d���roY�mH0��A)���3<3Vا����� �1\N�>�4��G��/Z'[�-I�s#��B�k�:P_nj�kll���eW���v{4L�q߸I���>�^A�{�e��?~�9��c	��89�a.;N�8��2o����h���k�����
"�K0���3# �����D����@w`� �@�[��O�R�R�Ik�l�z�n�SYd��w�ٴ��8�Q%�"��r�E"���ev��@'�ɕ��@���N��3�I��`�Fh�]���;��ޤc"D���" �]\<�=k�G$�Ť����x�n�-���k���nle�y�ٯ�)�@��q���] D(�
���v���u��+��N�B.7v�pr�E��r��^;z"̔�v�
�*P*�I;���->EB�3H9q�(}�*���ۨ�/=B����gc�V����[�k��Σ�dwS�6x�8�(��<5�֣��ge>9E?����e�p+/&R<��Š��(*���=- �OyW�T)�Z|�=F�������qg�^����\�����S���\���'rQ|�ta!#��J5����Fsx�K���h�K������Lp���x$v8�g���g+��sDwU@��}���}˕�k0"�j�_tV<��8� V�ǈ_�<`F�$n*�"����$r�-9�OY�����^WP�by1?���^�c/��>_���o�$*�ƈ;X�D5Z}�o�+C�֌���$��U��jP ޝPo���a��"��&�\���ｭuV�8�%�tN�WMLV�Vu)�wC�P�ӕtպ�O-'���Ds�'�A�ElLA��m�r<{�|��-��a�o��VFs�J`�?!��/1�c��R�Ѕ����f���d��$H���:���lf����+���!��?��6��~�Ol�a[��ݕ�+Ͷ��՚2U7���ઞ��/�57�=q��;SC�Sg��a;2JE�&@���V���{ц��|Amdr�N�uO���� J�
��f�i�u�Ʃ��&3��{��o@��IӤg�/��tP.� � (4jgJN��^	\<f�|O[�\�|n�ݖX��G l�0i��LZ�m��pL��ξ��ԟ��ǤR��>w2ڿPٺ�[��$��$ԸN�L�'�)�JA�A����vq5�m��_�]	M�%C�J���&��&Čo�Π��#�@�&�����C�����6����*��;���h���я{ZL.͏�`���5t؋�[��>]��0hi��+�������pV�L�a�ݬ�������" ���e��O@J�d�Ü[ߗi��;�g���z��w��I�Py���)�� ��٧N�ۜz���m����4������f�c:��M�����e�.���H�OD�>
�Ǹ5$Q�Z�l��A���B{�����.��gB%�a6g��'fޔ6���A����f�%j�X��H��C����fۏ��9���қ�1ww����0uʸ��Jb|0iM���+k������/�G�4I�ן�eS��x��� �a)j�r���
����+��i���ד����[wS���y���������FQ%��ػ�=�ޭ��k���9]��M*��*�f�^t�by��ll{@�h�<���\]�)A��0���jB58�vr7@��`:X�����ц���!.[���v�TѸM���aa46��2�r�&��mR?�3�~���^�i��Y�_��>��PEA�,�SN� Erf�[A��J�s�Sވ@���*��.i>�V84�����,�^�?�єG���k�Y��P�����9���Ck4���FuF�Q��E���vX#b?��T��ӱ�#h}�����y��	|����/�B�y8=��<�{;z��vU��o�B-���PO}=��KT����*���#Sx&	���"w���Ե�,�%N��7�\���北��5���D��zqq��G�ZE4Xo��9�|��	)y���d��F�/��6��\�����`�ե�-L��8���>�*���w��΍��;jfv�>�?]u�%g�0q�H6��-�y��cnW[H�������0և,���z·0������:�t4Z�Yt1~��?�P�Wp;b����v?z�Z�� &�4��r;hd����D�eO*f!�V���&�R�Ip=@u*I;5���?+}��+���l�ƥUz�:_A]I���]�6\�A�w������"c�{*8���)��T��ǳ��ަ�Jä���A�(�6Eu�N��6�u��"�m0L�N���*�yLD!���¼_��|l�\�O��V��h>xp�r�",��W�%���+�e5������?���ݛy�����m�l�Ag��Sⷹ�1�V�/;����+�Le�䲊��(��;W@�z�[TG7Q�%Pm��3�d���;�1�ۅ+�s϶e"G��&g0�/�M�����w��.|n�ǭ�a�8A�5�{�s.�cऌ��y�Ĳ��v��e��g��]��|��?�yW����F��E=h<���[����y�r�o���m΀EA�3J�B����$4�l�H6Y����ب!�ߚ-�p�%W��}N�����}�M��̧�����q���Kٰ��4a�����rc�o�N�,ʭs�������)Kqz\���tyi.
�R�)�ɮ0�Gp��?m�B���Q�&9�&�Cz�����r=kΐ::A��;�O@�Qd�Y��H-�a�(Qye;�T٪�j���v��g,��xۇH3�7���zJ����Ź�m�x��)h}�/veq�?�d;#M�\�M�5��sC+♗��R]�r�"�z�n�nI�@����RrN5M�Hvyg|��EV������X���z'���	�}�ޚ�l��е����X�2��ۙc���2z96�eA�p1|��Ǜ$�pI`��v�Vgg)Vle
+3����WԪ��sٸB$sd�NY7'&�Xe�XE&����h�4vZ�g�˯(�i-g���p4��q�ư�ܞ4�+޹��7D5,,h�΂#t�3�S>a+>Ն)��+����n߮%��Mv�~�rZ�_WS���w�Y�Dd�<�~�7���lq,��j�'�������=4�0����}_���"�a8��=*K��Z�$�p@=�p3q���"��sŸ�/D�R���ğ8�f`p�a^�B0�]�4z�N�%��㍊A����U˯��.oɜG$9�Z�>��а�z��,���9�qz��j�(�a �3�{����>�71����#H��p�~o:{��3����އ6�6��E H�KH�!�Z���(�*�$.�Y����ޚu��~������tC�x�Gst@��߸g��%�]��V����4՛���0���9OZR��:@���zb|��Nd����6���t�x�m��7�RKS��̯�Z^�]��{~�Q���6ן]������E�b?��:�eu�z\�{JrD��㮟�}��B�៖���b�:v��WFw�����R��*����_A�K�'�u�o�Sy��?�d��p�� ��;��K��1&�1D����#S<����;�N?)ݥȞ����cx�f�6)��x~����q��y�F��}lf����P]���QYx�ޝ����p>��}�)�a�AA���Awq�h���R���"�mb��񄚀?�x�m�-���O��UE��r=��u_>�i2{v�j5�s�_���W��i��m^�e�@��c"�������J|�����J\.O�x���m��f�㡤3AҦ�Բ3�F�eOL^��ٌ�$��\iVe�l\I��X{�-�+�}��������b� e�sR���&yt�5x�JQ��F��	J�-�� "+,��-e]�{T<������BX��u�/��j� ��Ya�&IT��`~�MH<h=/9b0��޼���{v�����i�&:VF��D��X���ee�w�4��V'��I6��~��x��	�s�~A�Ci�s̩��eT�M��$�22�[�צ�۞o�䨛����q�¸�!�P	q|�z�f- ��WZĢ���t�l�U�:��ӛ+��Q�E@z��n�0��Zl�C�5~]藮�t�g�d%.��s*��ݎ������u_/�O���4dB�M�R4�3T�	K�:�:}�^.P�S����&ޯ�(/�b|<~���H���y�q�V�i��n;Jb��'��!x��_��*���$�;��-����^5�$���1����;�
1��3m���d;�H��m�����"�eΓ�T����j�A�&Sl:U[[��b� ���U�flx,[v�Y�,�Ma�
 ��n_к	��c��u �T�/!�& �d׷&&������iO\\�;�#Q��	�g#��c���"/��F���}y������c��`�7D�ۧ�8O�b���{����s�NQO��7}�r�,������g��~����rU*�$��{�4�(�Y�$�ow�%��l�y�k �W�����=��יi�C;_c?Y:�6���~����H����ƚӁ��#��D��Ql���Mj��6�΢���G�\?��G���[�>8�ƥd��Mrm6[4R{N7��):��Q�{k�e	���l��3{��`�<Pi�<(㭗�o�`�-�`�Q��F�i����;Y���9�&Q�UO�C����d�akg� ���?u�#�pF����N�i�2���]h0�~�db�ja�a����3�:�I�Fx�H.��~�/�{��Nv>:S�?7�@��b�Z����o�9��&O50����ʮ�10N\ﺿZ�����Г���F;�u���ѣ��H
m��j�������m�3;�&Y#�D�?���8t��77|��wc��|�S��G%N���;��ٓS�pǓ����MZ�_oYU��W�>�+�v�oXW1�@:����{����"��D�U2��i�E�k�w���0�Č�X6�%m�� ֤��:�dB�*:;ei![��q�Ҋ���I�Y7V���i�m�;G˘FS��CО������%�3�,��R��<���	��3㰣���9z+��s��� a-��dfei˒����Do����iA�~+I�����t�����F6"r;��jq1�^y�mgX����;ѷ^w3��4-W��g���ff�U�N��f��z�Nŏ�Y��6���2f�Wn��!���{�1���WII�6���F8�3h�'Vp�X�)�˂b>���L��^J���c�|�}i�ͺ^��M���RD�0��oixԁ��T�:��d�r�{tc��B���PY��fz:�����T�<^����=��
u�����߼��F�����XWx���Yr�k��Us��t:�%�BaQu3����I��/�$MG4�G��J�8��[]���y�����E,��(Et���jE_��؎�����|�sif��¶j����IXd�����#��
D=����I�j��cg!X��]L��Ůx�8�-�"z���)?51]t��g�����ކ�񮻝?����WH��'Mh'�C����Хh�Ʊ.���쿘,�"�YF�%Ѥ80��GC�&ʵ�-eԳ�n�ڭ�.�-'�<�Q�����[GG���{�\OaH,��b`eȺs�J��E��#D�Ǥ��բ��4������iX�RB�����N�h9�)�)�ny�=�����wk�|����
�`@����(>�</�v���!��O7x�k-Y�y7�0�0�S�����2V�u�8���Mb�|�:�U]�렉9����fa;�x4S�I�,�@���n
�cxM� 2a���ef�/�U	����?�����_�?w�7�?��
nKp$ۖ�����O<մ�e�}ؑ�x��~˫W�M���@Ʀ�������.u�ƹ*�uv�;���r�8ظ����_ޭ�t{4]�Cs"�"��Z��"� �S��6���[E�<�����m�.$iZ�K}��a��39M7z������]�"r&��R'e=��ǟ��
����>�)�-d��d�ʮ��f��m��~lZlӼk:P��StT�^��ı�P*��zC�*�n��x��9���!Zx�D6e��.�^C��7t�P&Ӫ�����a=B�>�r�w�χ�`u��33�����,�D7{���?�	2x��9!����X�K��	�O�w��,��|�y@��ǦS�:rt�p>9�I.v��eJQev:��P��a?�E�V��9
��x�ݻ��=��iZW��1�)���}�W"1����'B�rp�E �������D��-�� ���З)
F!9�+�ɀ2)g���j�'2�3���Q��Ң��~ljk ��AS���v�y�89#�g�&=��U�y(l�c����W�>��i4����W%���RMN��S+?R�_
�E�
?ݗQ��j�V��D��/�	��]KW�����8pW ���3�f���~.��q�(Ļ�瑭��UU�6ȅ͸x��������������r��#�u�d!̃D�j7��+�G�`&����|i��x�ad{�~�y��D����}�v�nV��(�6��'��eb݌��3Sp�_h��؈��ny���u�Ʉ�x���<���t��5D���b�d��A9���:���qvz��6�1���i� BCދ����g�y�&�(�)"�A�4������2����>&�n޴��8��O�i���X����V�&�U�ؤ"�ګ����Ω�,!'.��N�'/$�Dn;h�2�D�q:��j$��j���u��;I�3[�����&�d����й!ҩ�V| fN�}°ݯX�J�%�L���3Ϳ�����
r���˛�D*������w�&-�H��L���kG;�
�]��v����H��� �] �56a1�.M��p�y��[?\}	.+�:X�*	�?93:L�0�^�bݜMn,�ӡ$:�Xn)V�-�=�bVA&XA�UƐ����
�x��qZ��i�j��M�=4���g{!1&��u��:&�J�KGv�`G
:�V�Π5՜��&�2��;Qx_�6��{;�j]�i]�-<�V$�5�u,#=��L;��}3��A���<���$�������-�YXb��ᮅ��+\sv���]z��G�)�$�?���Q�)P���9�
�\4^nlq7}t�㫧�����������:��c�Í�v�����FmY�a�+}�0��@C>�Y��y�!�]��>_οx&~�#����W<�`d���;=� �+QFLZY�����Y��R��X�pmvmc�D��tO][�Hx�W�d�����������h��(���3�
�w�ç���Ⱛ���q ��c5U���#�d�j�EC�@���3��as��}!�� R���x�i�Nq���V����$�!�'�mLZ�| u^3>���dIB�wo�&���Kd�ܐ��?��I���jD�*�j��#a4�M���T콟�G*���UϞ���܍z�ʯ�>%mL��m��.�{��F�͡��T������Q> ��L�:r�Eȃ�6C�t��e�^�g�}'����'^���t�K���M�m��v�X��tR9�4o����U�{��rT����Q����a�������1�+CWi*�
	��N�]"U�,�"#	�{UŸ�t��5��i�b��KQM�xzL��~�1�����Ԯ.�K��R�5���r˥��έtCu�e>��/)(
h�@s9����f�(E?�ޒE=�?����S�<�5�m�{9}�Z��X�g9h�e��9[���#G��|m�.H+�O3�F�u���y;�8��1��si(���=f���	}��Ӈt��Y��`��ȴ��0���˦3�L���A�Y)�� ���S�������6�iW����2�^�*3꫊O��ɞ�#��ӡJ��P1���/�.W���j�Z���6��X9[ ��v�bj.\/� J{�$�B�������1�=�����o�a���~��e�f�
��ɰ�4N!�g1j������̬ص����B��w��V��#Z��*s�1]Z#�ȱ�L�WϤ�8��A]�s��v��O<We���Y�W~gO׍�E?5ֈ	�3�5�m��?�������-�_��Pw2ao��t�@�'d��2����'3�=��d&�T���`o/��߼���\�'�,���?YBA��\�����+�Sr�$r?z ?Zj�&��0H)�(�rJ�?
Pף����5����es��|��w�)�)�x���7��V�^��o|�pf�N���|�~q��ҽ>�\��Sf�CH�S^6�SP]���I��:�hhE��2���ys̒����$����zЅ�{��U�d����h�=2��b�'b�vg���}н[ʏZ�������5\��w��O銆�1�>Tf��q�=�	TM{>/b�%F'���,�4��>�l3���4ߢ派jmd�lj!��Y���v�������0���8~�|1s�P�u�.c뚀��Ϫ����zd�3om���w	�a�v�&����\t�;2%������tz�b!�A���c5H>ffy/s�= ��Y�2�ir;��SI�=P���Ha��ve�\��S�n�7g��Ke�<FQδx)��s4�.?#(���9|�wH��=WnJ��[gp9�
�v5�9K<�`RSKQj�Aq�^�:�<��`�� �� �S�v"��[2#Ri"�Vl���J6;g��e��S+���K�ۿ?��)Lㆣ�\�㽋$���B�g��p��u:7':���&~�;Y/H�)�C�9�5)��3� �库v��D��� f����?+kb��G�,�d��L%gaP$��Od���:q�z�
���;C�r���y��C���.��S�J���m��F�9�Yr��2�����}�.�f8�TR�g���C�]+J�lxxf8)�iA�{��թR׈����k:���OFǷu���̡0�n�m�9D.H�*2�pȵ�ɗqP <Yf]��;;	�OA^�!�'���N�ch1�Xy�q�����:���62r'����u��G�m|�oc�����-T��C�i�r�@����哔�	�)���3v����x�؀/S����t���k��l�_���(�����j�ES�5.Ī+h�֦B/[�تV� �(���=����6E�_��������y�y�_�'�s^�u�ۨ����;5���պ�췜1�'��	P�/N�,ng&S���B�}�	���.8K�=/��|�6J�#z�=uJ�������T��#nϗi���n�v`�����4��SD�[Ya>p���c�/�U(b+q�W�p��!ɏM��{/���:��T�* tu�L��Į8ziF��
{�/Ӂ��~y�fv�"gO�>�En�At�/�ki���;� ������	��>�������!�ɢ�xƘ���p?[�qq|�ʷ�C&��-K쾀�J�m26�1^� �8zhxh#�]ؾ�	0)VR���o���x�� �B����~�X����r�F�,���E<�����\\��٥[`=�ך2北�oZF`��zy�c��$Л6��Ƴ��1�̋o6k.��"��6�;�a��O��ߧXn�$EV���r��^�ƙ������
a}SԬ=�Ɵ\1�Y�?e?ӳ�:��]��Vײ4�Vf'"��渽��ᖲi�v������w�p��ϭ��~���io��z���Fe���=%�LAJ���Q!<5�ۃ&�Ra[ïZ��_��
�Q��7�?�������[*�v�ç	E+po��}G�wN���h����~T��<���PtbEk�]~;-T�a�YkM�ũ�D;��,);�L��Ƨ�Ie�[Ͱa��� *��i�9þu���TNc;�����{�W�?��sU)��	�V���W�$Gy6ԋx��*�=L8�=�V��RJ�"�}� [ðt�&h"�
@�+������P��@z-��5W���{'�|<_�+.��=>N��]��X{G�}on�F�x	��a�p����ڠ �%�u_��}-���ه���9��b��^گ��Yb�)W~΂8|]����͡�>u�e��� �u��`�  �C�p8Sen�b7'q2%^Y`^�u�ܰ�;����]놹Vj���2,m�Pk�nc��Q}�Yi�{�'v؆��..^d���t����@�4�t'�������ŋ9���᭐�M��FL��R��/���BO�SL�Js!-�We�*�ݥ�YΥ����Nԃ8#g�P�����\��r�S3ѭ/������)a������=�i������+0NEP�}�����zχ'�vC�[p���\1�}�̄&ɼ�4;�-G�� 6i��o*�t��U����y��ԛ�qtl�!L����[.v����J�`���Ô���l���z/�P~^�\S � ��H7�2�����}G8��>����F[�9!�7�{��$?��ڥr���W�ހ�56����?{�����q�TZz&���R�|�� ��
O�F����Nl)Y��<��	=y���� :B8���m��n��8�����R�|6������C�g�e���y��lcq�x���v?���;<;��e������tE3M�!TtlR�t*��l��]9��r���U�MXu(�IzzcZ����NɍF7ww�Z ��«l�A1��r��dt�l+��@��R���l?1sH���?,~��qP|��A�k�B��j���{���@�Ht��K6�D㕟�
�3���K[N���T�?y�P�7�o g|���);W��L��=f⓵�Wc��z����j,���Y����y�� ��[�D�~����9�]£K��^�����K���U!�J9�C���C��s �E���P��J[yޟܔ��ւ�K����ƒ��Y���֏��+aYV��˗;3�ᩛB{P"�yӶՑC�Get�6݃ i�4E�o]���������u��]ݟ��s�ԗZrV�[����>�r�
��G�����MH��@���~��)���T*����s���u�m�g�sx-9Ki�ōL;s%L�3��r{Y�f}�������:����=��d�?��Jߕc�1�h- ����ݺ����	/�lGc�߀����,N�(�F������d��|�'�1���~�=�fc��>^4tf�V�����YT�;R�h�N~Ê2����;��?*o��
�;��^��\{k�u�����'�.�KK_;��m|�O��0�5�^�v,e�!HM�n�#�ng��Բ+,dQ.��a�]��qz,�%��`z���a	./C�dH�ţ
�H�B��z%hn����,f3==�rO<h�� )}pno샶�.�0ӕ�Spp?\��������S5ШC�g�f���I�;//��R�Buh�K$EC� �#;f��+�ާ����9[K��Y���;��l�1`Z(>��Lj=�n��X�;UV��/�M�Cٹ���W.^��د ��ُ�0;16v���	��¡Bj0��`[f4�5l��3������T؋ N�h�����a�N:]YM�����5J��@5c�n+r��Wr]K��E�_��#�
�n�=\�����+��mʇ��16�2�
��ә��� �	X�-Ɗ�PVȡ�<K�\���#4}�A�^-�%c������IԂ7�w�21c�*Y�}:T����)��wv�!��ph��m%^1ҏK.���(��w�`�}������U��zjH�?�����y�6F�)LfSט���[�����#Ż8^~%��f�nrȪĦ5��)�O����#�f�n]�uN�TT�٬�=/���M�{z�gmX�I��d�/��	�v����8���W{�7�����<&Aݥ�����i�k<�eK���ns���(u�-z$�l��R�9����O�����\�0Nv)���4��2)�C>��[@Ox�P%1�1��ܒ7��r�d�K}�﷖���%�H`��P}G�k�"�� �0�8�z�п��_�<��՜؞	��+m�S8X��P�S���导(�$�u>�J��W)t���U]�4oǚ밯���iC�(9ܒ�ll���}���9n��!c~Z��]��P�j���c�ڔ_��2���N@�Bd��^��ء93��=M�� �B�#��n�up�7����B��^�|�<W��6~{�E�p���UJ0���*�9$z-�d��&��9;X�aj�CN�9�+W��p�6���i#o���^��A�L�����x�F�9�Uz�+��r�oxL�A��I������^�(�{o���_S�⁏:gu����U3n]��M���|U�󹼚|�Is���mp<u@p+l6jo�ƠU��H�Ձ;j�o'�V_
y��ޛYW��3�P:�Ez�ڕ����T-�=Zm�LJ�7_����j�3�F9w��
J3i�� 8U�W@�81����gkX0�iF0؜�>?Bo�C�;��{�Qӗ����GF[K��	^V�'���jv���<�Jr����8$Q��Vf�8n�0��Nr�fr���*hUn��I�����1ԭl��G�2�n�q�kR��A��y�z&��=���6��LF!��H�?� �S�]�b���M��'Z7A]?���~�d{O�q�D��IQ�O��I�䌟�b�/jB���\bRN������tS�R�fI�PG��$��m�%M�<MqJ�@�ȭ/�ĵ�k�	*v��C]�-�]f��gۙo�Z��t��8c��SGX���}~*$e��W3:�iWqm��Z��p��+�����&��ɹ��g�)�O��Of�d�dm�XA��G7��n�կ	������6���_�F�o0Y����2��C���T�����i؂a����H�׺�Vg%��ڴ���;�	�wR�W�NMz�5�?�������`[%/���У~���z������gOV��8O�A-ͯ����T߲��PK   6}�X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   6}�X���]  [  /   images/cbec1558-c992-4de5-91c3-4ac90e5ffec0.png���S��i���S��>�����TJA� )��:��8I)�����Ox?�������~gؙ�$���@ �����#_>z' �1���<��K������������1I�n�g����q�~�����r��q�?�g�����VS1*8($Me�^]9�{ؐ���D7-;��ݣp����ԸT%�Q���%�B�ބqT��|>Z::o��x�A�4�3:߸�(ep�t����� ô�r���7�][7��G�ч���e��Ӭ��P����?�����dޏ�+3� ��O�W���U�����{���R0��Y��,��.����/ES�X��㺐��7���ZO���qlll_I�
XZY�ɩ�������/�?�?Dof 1�͏��>5U6w8��&(�l(�K��*�iyH��MU29��=�,���N�z|��;"��sQ�\BJ�<P�����kt�S"�*��ǘN�F,#�O}�T
kO��0?��s\�#������k(��u�д�F���]:���	׹b�w�)�5��b�r���D6x���NT�n�O��r�f��a���������JR�1m����СUPJ��1�6_��]���~Z���.����B2��Ŗ�
�S���Pp$q��%�O�k��[�ph%T�v<=9M#*����[2��}qA����h�!�0TT@���IC}o����	��� \Wv��v�霾�n��G����H���ե�ہ,2�D̍�Mhq�p�A�c�.P�~�ϛ�S	��E�F�,��J�:��@�EA�=��u@&�I�5���o�sg���J	���q`\y�#t+K��7��&8&�s8��$��ag�bY����L�:)p������m��9QG n>wU��	1cYNoqc�������'9����H�o�����(�:��_y��YS'��K��($H�XJ���Ox��\0Kr�DF�>J����z�?�7E�:�0������If��'S�6����Z��j�)��qZ(�>Tѻbz�_�J�K��sX��7vF�T��:P1������vf�C�a��+��,dK)�#���@�dy�\�ͫ2��zKB���\�,����2r�<�_u��^�U*�!��6ut-w5����e	L��)i�KG��I�L�r�S���`8?E� xaaV]����0���k�\&W������s�ؽ�*�-Y��U�=Z�����[��}�xOy����:/�P���r��s��+�w��׸�b�bm�F°�(�hj�l>b�S5��)���3��Oo��/?�?]e��F�_4T�R�0�}�u���{���iѱ�2=��CS���rLm�w��TA W��5^3�>����w���bܪ����%y"Mj\�2Zim������_�$�p������~�����~�:�������׉����w3(M;�ᬣ�L�GBҗVp�i�>�V�\.���e�êJ�/-{g�>8Z�w��E��O����ȴ��N$
��b��~���z����>P��לq�И*��L���ka��BƷ�'���̰1�W�)�у��#�|~B5w�5lX� �2�߬Bo8�s���h�I���ٳ�Dՙ#��?���:�Қ��+&�6y���hk�[�f�m�b��=f�� {�q� &�
ⱊ%�Ɋ��s���3���ט#�HA,��Ӛ���"�~�8�����#���q͞2Oz�Jg��`�"��*|\R���|dÙX�z���Q�Q6|��6��𱹻�����=�baf������������w�� Ip�8WB8���9��Th��ې�<*Z��/��' ɶ��7����d��� S�//Q��O��e�O���ā>y9+UJ!E�qg��:u�����5��{�������=Ҭ�Sd�l}*V���݄����aQ\���P��jO�+���3BѰ��:Y@����a�4c���ys�x���e���{ⲳ��n�mg�n#H�c��A��`�^X+����7KTVV���(O���熇�;�6^EB�1Gtaq�0J��m/�74+���%qF�6
�>Y,���ϟS���b P��O��D���H�;/ܗ766�m�p�L�a:�u/:*,$�%#���De����L9�a�M�ۓ������DTr���������z~>�s��͘.�[L�����͏�#�	nb�,i�3���7j����j.��v���5���WB�@��f�,��,rc!�?��αuZ�w]^9F5hC�444Έ���5���32��8Y�����S�l��[Q�d�ǽ������%� ��N������s��	�����21��33��#gg�CD^|�y&ʛ��E�:�e�����T��8;�K�;I3�IF�d�-gE�ao����z
a;}{rrrXUU�ܦ(��XFN��<=\ٙ�+�\��q���pR�{#&&��������&�M��� U�lv��όD"�!� �z@A�N��Y�j���_��^yz�>I:5�3�'[1b	�3fiJ��Wb1|�J=���gs|���"VK��II�p����w`[�ۍ"n�a�'�^s6����+�-rF��H��{���u:��d?�`6�l���$��`�O-5ޣ�w�LyÚ�t�e���ί_�����0?d� �n?ɦM�;~�}�T���-.����2'�z�Z��zS����%I#Z4[)���AR��-�j���z�/x^P�|�IR�Zg�5�ҏ��S�w�����Ӻ1@�V���D�JulM�z���>2Oo%LX+�IkЏ.��,��v[��0]vv�z�{$���P��_
�j�Z ��e��D���#�ͥj�oj�z/����6�$��n��܍p��4�D:g��'/�Ϙ��h�����f��[�We�\������N�+a�^�PӸBbXE ,D��*UPV�D} ���L2e���|�L�5:�Zjim��S��F�,F�E��w�B���0�ߨ����6�K���MS��:� �5�A�__�U!H�d��q�����1�M:��b]I�svVs����2}��a�7
;��y?�7�����n���Z/�Ifz��݁��/�*,5L��@n՛�"rT�[%��Q��}MpRG�����Qj�=1�=����'!��Zm��5���������!��U�>�#�5ߥ�(3}O��[�t80� a��P������-��Pd�����Q/��>O�\V�~��v���奦�W-u��5b��Z����1�i2�s�/_�P�����1	G��ks�"r��7�%s�jYL����_K�C��ɟk:l�����Ù��sP{����B��	xkJ{E�Vn�ί�_�4Q�/���/�uY���c�����cZa,ǅY�-��W&��]����*�n��Q})뵠�-+	���ڠ� �"SS���	+�"o�o��{G�ɛ���2*+�d릑�4�Y�ɍj����?KO`�Y�
���p�I���@��߄�gb����9|��wSp�?<��=�}�:��d��S9Փh±�Y�f�2S��ͧ��0�2�ܚN~�|W�I�2��b�PU�5�~��bm�F?�	-�V�zY��.\��U�S��veZ>��L�k�����������is��^��.���yz��t圕\�H0�3A,z�:~�Z�4�5*��Z��¥�������(;c�9�V&��"�Aq�TΠ�?��,e	��i���c�-��¹��*�x!F��Y\K��1�N�!���<�ۨ፩�6��4��'����K]Q>�<熉w��V=}��O<5��.ˈ}�}���y����b���Љꉌ�rdZ��.K�4�w[񧾿vf���pq�]@�e�me���3��޲G�zCBc��6�J=�|a3Ύ��$-��`9�w	��uT�0�����QaNMm0�H�5�[��DD'��s�!�����j0�6�ͫW;��YՋ��ͳ�ɂ
���a�7r���n~:Qفs�YU@�]�������#�o�$��/�Z3by.��R*��w־s����&QU���p8<
�S]GW��7j�Miˏ�-�/�:��?��Y&���*�R�̤�v?=;��В��	�JHHX�*ڍ5*�,j-��� n7������1��l&ۿD����Y�M����F�a�L�_��=$�K�b��Չ�}�n�z���O��E�@][��)�>�J����<;;$e���3.#���Al��ǿ�0���J�;$���:j%��'5h-�v ����<0	�4z>��e�r�A)]m�k4���[p�~{}Z |'>���#L�jll���W���%73�3����L�ޫ{YJ6~u��0�L�yq�(�,���r~�|4������Pͧ!�/��#�$XC�j
����o��(A��n`�ʳ��*
���&�?���Gs4]o�t9�	��zyOH�ˋ=��×j=��Bv���&��5�߭?�:	�� �� ���k���i�L�E}Vn�Y����ϗ?��'�Vo����{X"���BM�c4��(��L鐳�@����u1#>ǧ�Lm(�a)�RXۆ4�/�~S)�
Q��	@ӱK�ISe0�pj�?��;���fS}(�p�?����O��Nl꺲�ɟ�U���֮��6C���3�p�v�i��8�����p��)k˾�Iqc���O�	R�-�dy��k���!���T�tI1�LG�*�w��)z�]y
v�\s2<*��bA�IC�.Đ�����	n�!�wd{=����ϰt�E?�<R�w�_����pE�Oa�T� ��6]$r���^������)�~e:Y�&_� ϏH�,U:��`��@-�
���Fӭ�M*m�Z�X�Ž�I�4�C���b�P�AR����.�=����5��I� zÏ�=�"�	WNt�5�z�L$��Wn@�Ḽ��K�+]�_�"Ti�_-h2�
?��(�K��0�JG׮`�H�r����bGu�#�J�TJ|Ww��8\Wj9ͨ�~,I�b
c���M�Ƒýaxh$(�6ģ�|?"�l#ļ^�w�\CڞGpV^��X�~ۯ�	��.�);v��ZZ��(��ZH}O�y��[K��>S�垎%U�!t�,�PRjg�����#�pn3����\זM�H�"w�?��&nqt8��p��)��W���L�p���up-������t��	�ęշ���$�gP;i��C��u��w�OKn�S�W:k���~�4?#S-8<2 �֟\����Ӭ��=�D�>L�W��h�����@1�PK   �z�X��/F��  ��  /   images/d4cdd597-5d42-4626-88f7-26875eb62832.png ;@Ŀ�PNG

   IHDR   �  w   `�3�   	pHYs  �  ��+  �RIDATx��}��U����קd2)$@� �����T\�����b�����E,��P�� ���R$"���H�(� 	I������=��޼d2d&�̲^>a޼y����{�=�{α�o�oc�o����7������a�mlpL�X�h�2{���;��C����vuwT������M_r�G.3#�7���{r����S�ryJ:��l6���^:���4	�V%�;���+����_��W:�݇�xo��<^�̬Y�h͚5�������|�~t�Yg^~�Qx�����n�i�뮻��<����Ţy�G�iQ��8��>��J����EG}����z�U'�x�[c�[�0^xᅶK.��w/���S>t�G���_h~�c��ܹs�������2���$��r��U�VA$�ʕ+m>mg���=����}���a�4I�y�w�%�\�N8�����{  �"���ðx���Xx�]w-�߃/�˟�袋�ݒsߢ���/~����2�K�~�s睷��OAX�z�J�P:cӚ��3[M�eT��aX�:�Y�g��]�����y_Zh>��C�O���3�������y�{i�������ۿ��M��ַF�oB,�H�;�:����x͟����o^�/|�7�cKq�-B�?��>����[n���V�s�=ȶ]�
E�811�T�O�G�kS�=�����p���}��ߵ�#�M�_Yb��GWg�(֞w�9�����O[y�������%�a���i&�7����'���3�8�ܟ��'ߦ�<6;a������΃~~�y�O}����I�_���~�dSG�'�Q�t��~�_�۟�̙���t�9��KO<���7�p�?�V?�p���[�x��)8���8���E���i^s�5�~��o����1ڌc���W_�3>��;������~����W�d�!C��Ü�cvj��5Qlx�4�+Ez׻��'�x��k���eq��%�\�Cڂ�Gi�o��z���;�^���(0p�DI���QVL_��O�����f#�~`���8���{���ݱ�ڊW����5oGDF*���6zF�^W�"zz���6���S��<������k�|���?�����Rɣ�O���F+8��Htp&�f]�7,�~C�al�`�#�J柿��������AJ��S�d��XB��@N������<�0`"��R����@L����4m�1gΜ%�C�b}Bh�H��燿�c�l�6�(�_�hQ�����	��,�q�Y�����6�=���a%�f�����,�u(m��^k4�H��T��(�ʊb
����>�Z����~��G?N�q���o�Ή�MK,���Ot$Ću��j��q?&볟��������r�`y��~��w���[y ,�G����dR�_�@��,�I�:�@8I �bq����s�Y�r�i��}������?!4/��%N�f�)k(\����?8� ��9�y晃|����r�2j�h9a�t�qןq�)4oގ"B�@��⹖-?+�
i70mlݒEM	a$��d�w���ݎ>��c���_/ᏜH�a|�+_9��/���KNwB%��"�5A x�������κ�?�j�h)a<��s����{|���Z��+5�>��w�5�	b#�⍬�t�^���H@H���t��O��s��i3&�����4��$����L^��%K����vۭ5f��0.���?����B���j��ƺ%+b0Z�p��'�e2._���}�s�Y_����Q���_��'�l�$�h�����-3�[JW]}�	7�t��=�V�9E�w$���R�U)Z�`[)ל�j)a\y���$W_}��4	㩧����=�n���;f)ŴYG�)�3QA����}��ٳ��|��ߟ�{k���Yok�!o��④���Θ={6������6��ʛ�c$�����s��丆u��w���~���������`%&���"�E�'�x�Zqݖ��z�#|�p�χ��(�ٸ�b��9�ݬ�a�
�,�ŋ�e��`%o�scJ��\��w��ElOO���'''�Q�eaX��b��R܈^t�A��CصU���|;��ΫV��@<��cq�i�5[FO�����9waÆ�o!=1O7���''X�Cs�8�9s���gvn��V�X�GBo��Römѩ@�K�.ݱeץ�cƌr��`��6E�Y��&n�vp9@<��N��ݴz��Zu��^{mF��zk�D���\�r����n�k4����n���v�A	�ʳ���Y8�r�I�1���3Zu���y���	CɾM��L|D���I�ܻ����fx��&�fs�&+a ����m���B�44�u<I�8u"RxN&�����e����(��0h+�u����M���{����I<ĘDb$��y��f�ey���,:F�Di+G�y��l&�ɇ��,�Z5ZnK&hnِI�~ɢ�� ]C������G�\t8�@��c$��pQS(�b���dA��fc��|f�@�1"[[�4�AFK&�RQyE1��5���
����300H��J̈́*�O �	W�8��H�����?1<����Ds�K���2+-�}�hp����f�ϙ8��3o}c}����\=�붌0���Z�!#�-8�4���A�@8q�v�����^.��.gC���9���r��	�ɐ�$�0 =��,˥B�P�c�%�#�$
�h#��l�ha�p�+��P)�d�-�n���E��b�,�q,�cK/p�;OVrVK��q ���4�<�!�`n!��rU�pŃh'1�To�s&9��$�J����i�ò��G�iG���pY��J%l�ǜ�䵵A0�6���@�=��N�)�O���;;��B��){Z�D��g����9xUIIĕ���ʥ���N�9'��9ژt���D,�)r�J@:�E]
1�F�o ���c�Kϟo��_��;�h�5�6�`D3�T��{"�p�iӧ�?��:�5%�ϻa=�S�d��-�-�1�'@�mSM$.rȾ�����|;��|��fϞ]?��w]s���9q��xԑ�w�GN���;�8ꨣ*,\^p[�nV�8X�/��ne�F��D2�ň�Mx��t�mw�׾��2�����p���W�"	H[s`���[r Z�c���ğjU�=t�O��m7�U�t3��4>�K?vʩ���k�������~�/���}h���{�;��v?&�4+���=������7�y��@���ض#�H�8o:�pL6'W2Z�i���&k�*qpHM�G��_͋��,:v��W�.~����¯��7��v=�����8�?�o��Ƅq�㤎�5�/)�9L�n`?�tJ�D�����f�6)ul@rj�i;�/��8��aۺp�O�-�e�Ϋo�麅�v���+���/���1������ʆa�`�$u4p'�d�Ԣ�-�N�g2�|	��d���c��W	.b�h��~3�h�X��������q��_[�^��/ް�N;�:��!-�Gn�V����c`4ńZr�͇��)�dd������;�v�u?y�G?vƒ���g}�/�4o���Oc�������;bƮ�5�p�U�!�}$���%`�W�a�7w�r�/��r��xξw�}��]��/��?劯~��Oo��дz��L(��BVV�M<�8Fw+���	#����s���=������Ww���;��e��Ѭ*\��u;I8���u����%�`����1��m�}�{�\r޹�]��.�={�eW���oY������1�b���%~�@�*�?0&��1}C��'?��3>�i��?�J�6
,>v�����u�ǎ�N(����ئ�@���ͦ�~=I9��������0�/�����s�����Cl��L���PTA|�u0�ZEbu-�7%a4ڙ|�!�F�W,�0ů0�~��#�f��a��'�p��Sn���w.\x����ͯ��l֚l�)��?���%�.�a[0�:�rW�S'{M>��5y��?9s��#�Ng�V�Z��o~�۷^x�E�IE��
s��խ��shp�֪�1�6Y1��x'��~�����A����.��9p�8�1��JW�Y��c�r4��&�X�=�9F���Oj��s����s���=�<󌫘����ȡ�������<�OB���9��0��D���G�͜9s���5�;����n9s������)V3��M��F�_$DӼc3r]�b�i����}���p]�*����n{<��7�Xr�Fͮ�̥E#^7�n��[9ZKʌ%
�y�<O��bq�����M�z�u��l�o���F�VϘ��dN��m��ZB9E�1Ls�V�PEl�g��9�m��.L,@�nR�'��ko�w�̖��d�$Y��N��Y�2�2��);_�1Fw�01���Z�㴮�ũ���e˖e�I��~�'�R6��Ea�:�C��δS�7��sX�R)�OW�ߣ��[������3�<=�Ѓ�����a��0�D$�E�b�?�R�Bm��F��ߴ�%
UK��8����������k��RƧ>��k_��SN���SNy��]���o������D�*���Ȓ��0&��3�o��V��R��^uC����oe���対��Q�}�����NZ�ti��;�8nqk`j"�)s.I<�5�MǞm+[=6��e�qI�]�,tH�Q������E�_�S�Rؘ*oZ��0Y�S�_�٥���?w���y�G�������s�����b��re�` Ҕ�S��M�M�16��L.� �@nj&���d��"a跿}d��~��Z;�BVG#����Bt�i��p�����?�~�d|���G��bT�������1g�Li�500 �o�m���Z��e�]�p�%�Ă}cS��x�)���'�J��A��f�1T�WZk"������\�믿
�DU���@.{���HED5�u�*�EIh�������ъ�C�}��-�@�R���䮩�b�������A��
�a{{A��_
,&�䁠�	~?����z�>2�E�d�7e��IŜ���*��ۻV�%%�@���(��fh`܊봮p
�$/��v�$�K�'���Hg$ҟ1�j�ƍ���˚��(�0�p���5�؍��0WenL$�\���	�8��c4�1�S��jPK��~;Q�uO8�1�J���h����8���8~����`&�k�U�u�!�>�ĸ)R��c�j���)x=���uK��Vr���I1`";���̶'Al�oܦ���ٔ�k�o$z�By�ιNKJ�LF�h�WM���uG�Ҟg�>��0l�YՊ+�-���O"<�~=��U�o��#�h�Z^�>�c��Sa���cL�X�dQļ�-9�X�x���-�Veܵ� l�^����L���X��Y��Wl�h���s�d�+Y�¤s�� �N;�v2I�Os��78����
è%�d2�f����i{{�@+�;a¸������ř�>��<�(�j2Yq�o)te�\Τ�����~��ex`�6a\|��Z�j���^{�<<[���':����UW]u��>���o_�`��M��	�#�Xj;Ԩ=��pR�@d󛬣ӦN�J���B8�?����p��_�c�׹�;N`>�T$?��{<��*�-�܃|{��C���#���?���i��0C	���8�t&�/7��,�>Dzz�!�7�8�+��leSn�H�:a��$��$:���P(��Ƅ	�Z��(�b�{'�K��
�o�N o8�Ht��cpp�mS��Nr:'�� �JUBMz^�D��&`C�rH�q�R�\.	xk�4@�X��k�x���r�f�Y�(�[�2I��V��'LȎ0:�<��@:)�R�,S�M@�^_�]�1i��Ġ�F��[�ӗFI&%�L�HI��tOE��e���D�1h��1�@�J������iH�#Al ]g$����0��O�t�ϲ�U�'��1,��@L�EO�\�%����	�sM����w7����,@ {ǟ�ST�BJ���}J��3?�,N�s������HH����wS9�����\�s�ąw�YoX���&�a����&?K����D���g����#���)ND?�*�)Su��b�'�3��L�;�ǡW�S����:H���xA�`�a}B��'L�m�N�u�������2i2� ��g��d6�c��	�f�!ʘ)�{ȟ�MaP�Uf��R�n���ɷl�XS�w.��_�f�đ"�Q8F�"z,e��'�I�Q(VM����G����uV��V�R|6Bз
���xD)��a��cC��M��Z���.�X�0�`���Pd?�C��a�:���EB�O�0�8�>����l~J*��j�Sh��3x�[)?��v�ƺ��N	�gx�"^�J�L�c�x`��0�+�O\��:,�׷�I�*Lm��̘�*��e&�����:>�`̵����Z1��e��aa`x�n��i�j���<0$��P��q�S�x�@��d���ab�ۓW�2��	�e�vT�Lc�p�g�͟*g̺�W�L�$�0a\�݋�����|�s)'���Z���d���~z������_�P�^ه�"k!4�����e�[��^`���:`�[5��&ˈ�}�&Fd�S����a��hC�D�k9�m��n�F�U��2�D��,�4��BoQ�^����C_���ڔ�|���O��''c�3V�Cx�s�]{-}����ț+�`����\8���+�h=����++���������|����Ь^�����+_U�}&5^��yU�_8�4�1a�8���y|�������rՊ���N�M}���'?��<�����[�CF�Ȼ�������p/M��5cƋ/�Y]�-E:��(���ul���,5$7cF[��[4���#�X�ݫ�Z�:��k>1����V�~Xd!Ϝ!8��&Q`T*7�s*�T'����a8�N[:AնxU�-vg�R���g	1�ޠ9'��y�rW�^K�Лc��k���J�8�2���yQ*��avEp[~���o��Lyh��2�N+��]��SO>��1���ʹ"/m�N:��N��u���o���z#������&<�|⫞�5��a6���i���cPkPF�[�0l;��e�2�Y���E����~߈�]���Ӱ��(2*�遨�S,v��I��������l�a�2���A4�e�6&[6�Ҵgm�1�0n��?�;�����:u�df���%N��<6��5����AZe�������wڐ�E5��c*�����Yfª8*6�{�:n"#e�3FD���15�f��K���Ղm
�TM}������B���H%Ū�;N��xm�>V�q<�Ib��f�v=2~z��~��j�H{��^s��7�ڊ�������]uH͇�{vY��ӴE^Y<Ł�=�Rۜ ��+�� �5n�7z�7F��l�1�]z�7?������O#�/N��q[��'��s3��&��1���t�)�GFF�����(ӂɏQǣ�l����:r���L;��^s��6yٖ�ڎ���sh��������>Y��Q��m�o��T(l�m�{��]�2�,�a�ෞ�e���J`K�cID7
׍!P뇬��\ެ�N����j��/��y�5p4��>�v=��΁0GE�c�v�1-�@����۳���(�e��ݨ�{�r�Ƌ<�۴׉;0��]��H!��M{6	,����
�A�ӑ����y�в!�R�y
����:'�`k�0e�qVN�6��z8���1���9�C�
a](d�Q�Lo�V*9��08p$3Q��4����<~�i��R���*Q���M�ԫ�O�;�����l+�E��0����5>-q�����.��h�.;�`��`e�ژ[�\�VU�{��S��R�����G$�v�ܝ2�IAy��R/Q���Y�y����e�yU�8�E�De��jmE�&F.\��ڱ���pb'O|�뼉v��7�9���Z��z��[��$�a	�p���K+�Ӯs����p�������P�_O��/�ܗ�A�]Z��E��TIt6�l��l��LhU������������p㭉������yÝ�M%6��TF����ub�H��z�H5w6Kܜx8�z������,����A}�=�LEU*�j��6�9M�"�?���akǕ.�&��}l(�APhR/�G�bA��iȿR�'�=��I�=���UQ�$�A⼍A�!��x�^�F�+ejgkg��D�gH&?�K�O��(*Ih��>?�_���PY�V��o�� N]lɬ��aȵ���R��<d��L�� ������FיS֘`�8>��e
m����2��^�~�}y�u�oh�,�01��L�Q*����ג��S?�bŘC��f�cJ�0���Iq�d�m�R�F��ވ�e���(�����"�%?m���]B�(G :�	�4��g�-O�R?�%B�� �hC�7��,�l҈=F���ұ@�G�
�#0a�g�̚󹙔�����	i�0�6"��X��ux��������ƈ�2F��U=1�R��O]v̧Y�P�;�?�A�d]b5مN&��{;��NN6Es+K�PVd�V��m�_��=�}�T	ҁ\+`�� b6�z����� .'��  T?+=�g�������r)
�a&eD�j��`q�C��D���qX��+�Y`�e�XD8F�O�"-��wl�~Z�6D�2�E��&/�̈́P���N�ya��!6f:�(��Ї�7̒�`H(*�f�XBw- �d�� L�ejc%���b��/%<^�E�����KT��M7vRi96�P����ׂ�����%�ʴ��R�t
�R�qP.�F�؇�7�y&e�GT4�� JF �G�����`����+��,X4~�]���l�͗0M��K�h�&�v��)�����x��L*��>X4C�
;)�^#r�<_���o?��h`�� AVȊZ�#VH����5h"����w"�G�χK�]�Akʒ�p�y,F|�T,f�>��1���+zP�D�C�d��"�L� ���L���X;,ZB_�"�!�m���3��I��2�tA��D�
0�V�b��9EԄA25GQ8sɄ�BJG�� ��e�?�)�J�]�����X"�J��|QF-��.�j���0D$�S>/�
>�7d!Գ(U�l,�0�J�r@��<bšDgRt3�����q�r�M�F�T����[�S��V��;�&%n���6���Ĉ���G��^4yc�Ԉ��6�$���(�6-�\H'�p��P�
�MWēMUb ����WFT$��m=m6>D_/䟞(%���D�Hq9C�|%>#э�rMj��P�91�y���#���{C�Ew
c��"�_���ޘ��|���3R8E�(�.�Cs:\_�|Yej��cXcG
3�5�Dk��^djq����;�R%��0�ݑ(�"!��9��P���'�D�C��W�/�J_��{$�(9���,�G$,�l&�	W?T�b�sX��
y�9e�B�
�iQB��}�ܲ��`��1��Q}O��8�|���(�0�c�F��(W��:5�Zdَbq��WT�v�T}�g��}@/*`G�՛Ĳ4ʊ��Uiu�;p��5C�e��D�	X�����	&��(9��f��p�^�H+�X�HqAc��J��4��v��H�[�8�1��>�d�����G�m�,�S�u'�>b�����BP�q}�R�5SDф�|V���x�.j�#6�M-�#q�Í��F��5�U�]�+�M�/L&(1g�������������X�bs.L)	����(�b7�[�2��B�ն�;��w�S$�Ѱ��~�h�T�,��<�Ta�_�
�{SX����8 n~����7#�,d(�4�h�4ŬS;
[�����xN3���"�E��j�ǉ�9�a��8Ƹn�(pvf��7�T�b���Q�Y�ld)U�PրUi�Y���bd�1��8���x��q�k(=A�%W�.N�9@鸇��6��6�H�~"1_�=\���&�и6a@y��3�\l��&��GyT%42��`�q0ڢ!�`]�b�ITi��xp�0O%�n��[X��Ӵ�G8m�1��q��NciKqb����	c\#VR���@�66��g�����O�� ea�D�(d��q�dL�K�&����/>���b�6s��J�T��UWe #��w�*�v�4d�4e%4N�F��L	���XU뺎��*:1�� g���i�h�9Hy��sfQ��$`�cS��aJ<@�a�邖���%bK�h�ڃ5��5��X�-�s�����#�g�Y�0aq7�{&0 I6N�8�bļ�,Y �f�E�B৞�z�Q��t�OJ�Mg�Ao`����Y��<�ê� ���������Ar��^��!�� ��'mJ����2q���sT�2�@��K����(�-��9�	,,�D��4k�:�<�2�4��I��< �: 8sr���T3�;�c����fnQ���i�[}�e����"B�j���w�b��mJ,V=;�&{�Z�Mִ�@F8�R=�aċ��J�.S�]y~�6f�i������W'7��)S�O��DQ���m�PDQ���xd;���xK��d��A?�d�����+N$J_�(Fù���P��fã;�!q!'��������H�O�Kވ��"T=�JL����
|_&p+�'+,�����aQY��?��3���+�e��,X���O4�ﻶ8�&:�h�$��W�'ɤ���9�M�ޫ�rh�e�c�H��H$�XIq�b#��0qYQo LS+ ߫0����+�H�Xs'^�����e�\Wi9��i���I�E���$M��	8�T�8���F��� �jHWg��Qۜ�C���"��:�ق�Ļ�(mz���ɅŐ%J9��L��e+/0�ϊ<b����	�X(s�1R�g���$FICX1���@�c��,�W���=}T(��*�F�
��,o��� �j�)�0��1�ɫiժ�|BJb� �������R���7�o��Z{� �IT���$�u!6I���Sy�^[��A4��K��1qx�:�9C/K��	ϟbQ�fh�LY�2_�.��:�N���(�#�f�N3����>�Hq�!Kt�(gieSG*C�ę���@,�b�����,�"�&�cK��F����UQe��㇅�Jj-���;�#�Y����W(�1A�9*ȸ)����;h(J�uR��X_�q����wS;�D�h$!oڀs*`�XW�5����l����O��sur&���Rm4�{��,�||��2hwQ��x>X�j��!�'�A��J�T*�y&�
�_�bT�c6�� J��1�'Fb�Xm�#*� /@�����4C^,�x9,V:�[%yRBA��X����	��Z�,k�a�5r�a����]1a���ڌ�tl'A<���iPܘ��}��t"Oղi0.(���q���!$y�E&�
s7q剗��P�]��\�N�_�����N��>d��C�X�*���� �o��&�Ԭ=���YN�<v�I"ǋ�:ZL.�j7j��m1�P��7S�6�S���r9��g&d���Krt�z�-`B>M��i����/1q�
��f��9֮s�Q�aa��FcP�L�����s<ǩ"&�&]�V�C�R3i��Aui�w��$��_�TYl�G�%L��c�e�N�)����}�,> �)��0��z!RO��56QbF�V@��i�1'OE֜ײ������s���ryuX��]_��ꄋ���^���*�;�l۲��>E=QAN[��XD �v����(�ǒ9��9��N	H�CQJ��<���F���	Ew	"�1aDl��R���Y�xc#�Zz�.�]L�Y����{2W�dR��fѐ�c������k�#�ֳh�W��Úc��G��D�&쨋��h=ǈt��j��)��Yc��'ކYa��~����L�U���@S��.3G���8iz%��o�	Wx+QM�O�9��Ma�s! }"�P���	#�,[��\
�T��"�Ֆ���32$Fo����x7S:��f"B#��b���u��>�F�:EA�0 ��u� )����(����U�_N�oX�QJ+��j=d��#��ۈ*�ߘ��U51��ŏ���2J�K�������ʬj��M�I�\�I���F .���zVEW��H]�H�F1��]��j�Ni��u�GM!�
b�/	T�U棸J,
ewF�x/Ԡg�pr�MQ�~���§��8u�W>�H=h(1I�B2��b�a�U�C!���0�8��L��= L=��5��&J�5��G	�N���t�ر������2���c
�K��]�K%)����^���rRH.S�bI��aE�"��Dj�L|�����Ig�ћ$M"V�6��� 55Ľ�Xob<B���3�1�B�u��g�5R�	_j��G#3���&!*xK��c�J4�h����$�@�{_��u���RJD�<�OLlDԌAR�K�B��j#"Smr�)4~.�HGx�i�@L�d�k�i����e����hXE�Òg�@#��"3�֐�`���¶N۰5��z�T>73�HF�s$�������J94����������a�a�cWU�� CgV�-�G�hK����6�c��9'��ǖ�M𼂫h�7�Ok�(C�.�M�Ex�r�)`��TF�4D!A���Ñ2UVL���%�BHEmC�)�J$vMPǰ���ݫج��vA`�á"- Ԃ�fɡV��u�-Pe>�B�x�n.�xf��@e�+(P�;��fJ`"B*��RJ���R�l�&z���@����:J�]�~}E4��E�w��|&U�-��s�Ɏ96D۬�$6��]�la�n��%2U��V��g�d��H��,Ca.BC��f�'p���@R��Vk5�]^ac�K�/�7��4C��" �%b�R1QD.��&���r=��|�8#�l��gR>[sE�Fl���:�9��G�ceu�C�� b-zH�*F���'��6	�3��6��uٮ���H>����QO����OB�tq�H@>��T|�]b�=��Q�[��K	�R���~C�Vt�0)3I�Y���ua+.c4�9��G��H/�Dt$�*��<�5	?�!bn���5��'�X�0�cC�������_]��U]JB��Pu*��'�~�ծ�C���C%*2���i�s�CQ�Ė��W of
KV-Q\-����g��p��@��P5�ee��بD#h`*c��K��Td�P"I<��b��\���馩ce(���U��YA��6�Y�9Y������r�� ��^�\�@�rI�c]Х�����t���|��m�i�	�75�GV<"�m��)R#3�K�xQw�;�-��������L�Hsg̢:9�3R�R�����ry�"��T;��p'^NW)���i�c�!{���w��uk������U��Ux�r�i�P7��c�)��ԙs9)�x��ixs��>�r�5��|�,���bţ0�Pn.[ ��VA
e�Y�dޥ��\�t�]\�N&+DЖM���NTJdY���Di�ζv���g�à��6�_ˇ���*���`�*�%�I�����ja�	cc�.I�x�b�Lg|?z�e�'�7P
������Y9{�fP��3�|ǟ��/�P��)���R�r�H��}팝��K3�6+ǚŮ���]������3�U�pTS�\*נx����R.��b�`�S:;��,xa8|��^@պ'Չ�s�Z�*��(�L�" �2b�gsm�;��5R���4���V���LA���v*R.D晋Ʈ4P*Q���JuO�7��2�<g�#�B*b��զ&��h=�����% `�o�#́�/jh.��57<G�y�L~o��3��3OڃY:@�W=A5�sYތH�Oc�&��A����e�Sɢ�5͞Ӭ��i��i4��#�u��D��5��L�u��a�`������6�������I�:�;�8T��y��������=��C]S
⓱b��������S-ɯ�T��ďA�j�ژ�Qq-�S̩�}�N>VS��w����+��)�E�P�Z�klvQҌ��U���T(�,>P�J�b�O@%v�hM�F��<
m�=����]��󎦽:��������Oh�L�����f*�]s�3��&N���g�C���V3[�@�4�4E�_�5����7���1�{��Ī�ۦS�u�����wҒ����;�F�z����^�ǖ,�߬�:+�(�]G@�Jo{�|�6�[�R���2�˫=��s���A����6��޵�n4�};Z��rzt�2ZSdn6c��F:�s�Ϗ>H��:�FE#Cw?��E^A��b�*9�/eM���;�=�@��	c>�2��$�2LV���cy�tC˱� wb�O5!Y�ev�V��%ϧ.6W�t,q���{�dyfO�z����TH���נR��U����B�$z�L��^��v���o{����_,"�0��2��3��ϡ}�a�Δ��Υ��w.�{�誟�KSXtt�N�s�NL5W�m>辍n[���0K�t�>�h�;�q��4�Ŝ飴]t�r���%T��m;��>w�,�ޟK'��?���h{�]�ɺ��}�mM�DԢ��K��C�jLS�X�o��u1�sR��xuCխ�ݩ��P����Þ����O=K�f�@eF
��TDَ<�q�+��_�N�6�˶���n�1+��n�~��(CCk_�?s<��D��@O/]EUՍ?L;���^T��*Ma֎�co�=EG��m������S[@�ٓ���K�����N#�+g|���O'��jƌ<�Ȁf���`G�&�Ǘ�x��.Ru���}���鵥���DN�j��D�ͫ�D�|��5�)�1���'&�%��8Nb��T�e6��gd�c�Cec'�J��.E�L�WV��j��rJU�>�߼�������މ���V��T���Ot�^�U+ג��A��p31�����=����)8��t��t����>���|���_)�wSG[��Ţg]A/��Y*t�(Up������Bއ����Rɤ���G��ȓ�ߖ�~�`���=w������~�`0my�ӦvRƝFC3�r]�T+�N:R�q��p;���g�a���.��t��С{̡�|��W6�7����>�gr;w��U@�6[=�H$Ш�P�D_Z^e���h����H<��M���T���c&c�-rT_��,>}#���K'���t���oK����CV�2)��E�jm�X"��&�,��;�?��~������_!�}Gr]��̻aV�	�urbjZ�n��g��wn5h�C���}|;�cv�~��g�}j�fg���:���O� /��"Ųf��X`���=g������&������W���<��{������˾y
=�2s�_<NO=��ܮn��Y9�E��{eo?��S%9{���K˗	G�u�)R��ηK��g_x���v&��L�
�$�}�e�R�*	��;Q�vC�j�nc�4GUhA����C<�JG�y�$�ꬿ1�Jƍ���Nk�B��O��=_��6Ņ�*��zY�ɰY����>�	H������}����NL�_�yz�Q�Ko���A��LA�TI�R��葕颊��H�m����u}�����L�;�$č�zm�z�dQ�Γ_���ZCKW������f�B\b��������VV�}�ܛh���л�K��>��g���C=���)}}��Nz�C�C},��R��M�*���YJg34X,��`�:��"+�[gp�	�(�E�P�W�!�C�FO��=�Di�����,�H�(���[_i�[@���]�3R���VO�
�%��03���̲1i�tɝ:�V+���W�>���nt����1�?�[j�兒�5Xe��k�f��YNէ뮿��z�I4�Z��2)F��*��7�G~��t�G����ffS-T�.L�[W&�Jp���8)�'�*�*�f3a9y���ӭ�Wҭ����oٖ.:k�y��韮�9��uLgQӖ�� �M݆*}EVZۉi� @�V�؄-I�:9<�+�XgE<�fn���W��Т[��ſj8B$k�u�*cH삂��m)���@"k,e������g!,��_<a*�'��)��&"nqKN��e%U1���z�CA�ewz:���􁃷�SNؙ~��+R�=9�٬@�C��U�y����֮RT��>�@��˯��5��5D{�-��c��S{�@��O�7{6E�L9�(Y)��&��,[E�j/�Cm�5[(��@Zߚ54���?��O=F=����N�V3Kx�W��mK��so�颧�(W���#=PD�ݿ{�RLxq�� /W���1��L$�C>����pB1�"��L����R�0��4
.j�b��0b�{A���oF�['�W"8�並�*�@$�t2L �����L�G�Iz�C��R���H����|�?[����˶��7<E�|��t�GХW�GS�fP=����Ot�ns�c����DԻf�,����=w1��'�0�X�L�MW��t������s��ޗ�^�mfmO;��AW^�$�i�R>}3�d�Q-����T��9�O���Y;����h�w��I䱂�ڒ?S�����hG�W��˄m�ѿ�F��mK��z˜����>Ms�sz�M�����WXL�ie����X� bf��0'AV�ҋ�fPcˌ���d$Y=*4���*a�t<%��a��.�k)�16s5�6ݏ�S����$)EGU��zN�i� ѫ��t2�~z
=����f��LTO�iy碷�n��l.�؆�eJ�w�@�����
�|�4�f�c[*��'���_��=�2��N�ryz�%t��K���^:�sD4�ġ��Ѳ���A��
���Y})��ζ.�f���f���c��N9r�cޮ��S�_K�_��D����,�"Χ�^r}����C����'�f�r��k��w>Jv���c�;OO� Zœ�����S�4"�ď�RcV����ƪ4�I&���^(d�ш�*���!�	����F�%E	�3�S����.��`
T�M��s�J6���`��ѓ���w/b{{;�U�6���x�T������28eZ7[Lrn���֣~���L������`����g��B��V�C�C����=�)���W�be�����P��K��U�εI���`���^���>��{�k�j�nz`�tσ��D��NQ�Q��]X5�K��k��ϟ��n7���*��<�X2 �e����^��K^�+���ɢ�g_�;R ��JRyQx�(��.����+�N2O�hbH��e������p�&����g�~A�L���� �����S�PQWVP���uH�j�/	�>@	Hf��w���Q�!h�Fqp�P��FTc�5t;�$!��i�WA
CPS����)TD�8+���`_ޜ���b�L��,6��J	'B�ӻ����_���i;�[G���HY�q2�C�mn�#P��$�XJO�#��k,G>����p�Ä���!��ܬ�d �{K��b�l��3V����4x(�b�O���aB��Gg�t����@��q�p��o�v/�k"�
�S���ME9�5/}_`.���B��À	�C�'9]"�,S����P�[ .*�,-m
���*�WbK()m���A�=�m�+b�s��B`{��Ҩ�㤔R͛�+�F�g?	3�����������
Ѻ��<�X�%��B(=���ʉba�l�j�l]��a����*.p�=c���Y�'&VR�-䚘�n�
,���_�V�RA�H}2�GUAccI Nc!��U��G�e��J@��7�AJ?M�O�@���T=T�A��T
EN|i!)�Qc��P7(.����Cĕ)�{2�Ȗ������n��Mq/��#�%a��s1���"���b��(�^�RU��������� ��!PB�-��,Sk�MJ��!�rb�5' ��p�T�J����Zj����G�A[���yҗ�?���QT�ut5�WY|�'�<��/�k;��0�y1@��U�S���wL��NDo9a[�п��yA�@��*a9�eE�/R��Q����X�6�t"g�)Ś���V��/�`��'R�l$ʲI�Y^ &D�!@8 Ѡ{uʲ�$ռX
Jy���l��5\�y���8�R@N��8�9(Ub��3�V����0��t�s�
��d�mR����8�XԘn�P��V��51E�Y�x�� ��͵���<�����T
]Ή��pe]��]pٔ�P�֕ �X<�K���<���(
�b���yUI�����C� 5��U���	`�+tba��	��v�R�+��,��eQ���	��h��I��@�����ErA�<�j��rA<ӑT��-&$p+�l�.��M: �D.��1� ���LmF�C���!��݉�`���	��@8�ͬޯ�s�r��t@2T��@O��a�5 �
O�*�T����e3қb�R~X1��@2oul��\>��t#I�,y�A��٬bV�PJ���׵�(��6{FG�8Y9ˣ�W�P��*�_���f҂R
�jC�h� ����8�N�ιT���IʋfI�;X�S`�Pz�E�{��L&(xUQ|%��*W� !@�\p� �w6!�)����s1,0�[&B�yl+�,����Tx��[$Y�!0���y}͛
L)����!g�n������,:@U�O�*}+�//�bsHǄ��e̛��k�G���*��<Wg:M�>�� R����gB˸!�X'q��4��%�mTS�@w|B�^�s]�H}Op|��v�ڶ��(�Tc=��=��1J��1���U#��+7^I�Dk���$`(]@C��A$�
�w4��mw��Ա��T\�Q�*$������釩��Ս�0�+T�.��U�V�-�l!̢]�؎��4Q! .^�s��O�-�5��x?��TH�*u�G���z�#s�&;�N����̳V�����]�C/>��'���ST�~K圲|ϰ�8F5u}��#p�}h��?C%t(w��D�c"��x���??I�������v�K���!uN��5P��/���?w!��n�i�������A�o���@���g~��e�����(�0XT��-�4��L&G�����IauP���l�y�!�A�'�v�9��y���
��{���B��N�QřT�'�レW������_,�c����\CJ&�L�Pl��#^�iوf�;�v�1�Y�R��k��9�)���Eǭ��AO,롔W!�S��<s�|�u���\L��wo:e���5m�A�ʞ�,��3Xl�T�n��b���s��l���e��0���Ru�������fNTa�H�/b��h�DA.27~�5t�od�X�����'}�bS�3"~�'��1�5�E��\���6D�n,09'@[&պ
� �D4��giv;��� �Ѽ�	�w�芹�O!��Q[.m�������󑥓yP#�9�\�)Lp]i���*���7|D)E�;�i�	������+�E��iR��Y�E
���H~2���x���# i*�ZET{����M{��Ւ������b���b��כ��� n���q!��q�c�YA.�/�k���^#�Q#ҡt�cBj��F���*K��|�����pC�Ft���kؔ�H꧅��}��iC�e�uO��@�fٌ�E�2��{6��rq���4���3a��|���AJB�p �ԅ�&f�_3���&I���9�p�C�ur"#V�Z�� rB���$B�H�M�	���TX������%׍'u�F=P�bCu0lG5�&�R�R�M�+����q��|�8Pu� f��bԓ����F!:D��y�9N�)����
U44�k���5���yD��bh��-�_��÷�z��Q���~ �lE�ե�)C&�H7��m 6���cH G��(�v��L���-~~P$��R�����n�@��sǺ�f$VNzv�=���4t���2Y�W ��#
!kZ�����bV��L�)1W�r�4BK����gJ��##����瘽{��=� _��-���T�3y$���`H?�x�j]�d�\Z���J<��T�*�L�_I���t.��1p�2��=ߴ.�y����etKJ���{�:�M�Yʁ��߈Ԏ	<ޤf&�� l�*���}�ڵ�7����F��]�d@6By��,�8#�k8�$0��,�\I�'�(p�pU�$����K�Z�|���Hm8E)J�d�Rg�@�#I@B<:���T�"!vd���ä��@�Ռ���
C����J ��b*M�:��T�@E��GWrz-d��򘉠�x�̭`���)I 5?���Q�IٮqA��[8�Ⰱw�y'-^t�,8F6�j�~��E����˧�$�9m]$o��p�.^�.���
���:f ��iB�C�It���ZU�P`�H�_��T𹧞x�.|�/��N�J��}dQxA+v�WgQ�1�\ fE� .��"�^��sK�H�ܼ��H&rTsa$U�	�b
��z��]Ya1���Ɛ1\�UED#���(�?��ZJ�C��tEUX>lt�d��M��\P³&Y�9o�����5��%�!<�._Nk�RcS���q�r͆	
�){���]��c7Q�g��Q����^~��[Ջ��\%��~�4.��F,7|��R!2��¢�� �4ܲe�؊,�e��9� �NA�����i�+�C�T�PA�j|(�lGC�����ء����]R0=f��w��(��দ����a��Ǥ�[�,��T�$�Wzı���֧�s(�h�ƕ{`�c�ch}e�S���/7���C÷�:�&i!jd#`%�I}��l"�憱�!l|����7��-uC��b�I)�O)g���M��i�?��u95�>r�x��-�v7gش���t�q�aȦ&!p)0N� 7 ��=G7߷f8�~�ah�/8�'�8���~U��P}\��bC��J`Ѫ�}t��h]
i��n�f6,�&|�F�HQ2�lwY�jU60�\uBI���.RM[�H��}�D̤R���e��ͷO^�̵f�1��IZ����{:�3Ho�с>(���@�MD�noXA��'=�M�8<GC+¢�e�&�,4�Q��U,�()����d�|H��@�tD�F&Y�h���EJƽ./)nR)P��zS:Gi���T���b���+�F�
$��G%"{�j5N�p�X�G�ԼF^/f�����hː,r�g$'�AZ�l���=4T_5�u'�l���9�b%�ћ,�cP��O��zC)��q��M�Xx-�H��b��*�I\+�8,5��~*��V�VR�]B�Y�YI4�~����'8ҏ�DY�.����DJ���N=���L��Xz$l]m*563�UJ���aqE��d��6�q�Z��78�*����5�&�����Ł�:�(D��'�o�������:����A(�X��$��֩���br;�5G��i�u�HS�DFb�V�+)�I!�ULE\|r�tbQ�j�XR�Η�R��A���]R����|n�\�kl�jQ� wx�MK��_���F�"��Hİ�qZ�L]K'V�U~���|�:���0��Oƨ�����olA��S�E�tm��X�%f2D�IM�XNw�X���0�D�$AB�����7)
&iAb͑٤�5�X�r�H�q�J�׎�EL#=.ɻj��O<��-BE�5�'�
bڊ�%��F����b��0�M��#H8���/z2�eS�8N乮5ּß3�T��M;���Z8ĉ&@�@b�(����Nn�7^b=ڿ�|�GҬ���$��\�x	Qp������Es&���Yqn�|�5"�r�?#J��@�,�z[��@�Z
*a(΀^1D|F{mEq�_ƺy!� Z�|����4�Q��x��{��ـ��3}M�\�ډ���xƖԝ�8@�eDB�]�E��<)&�>�&�$Wץt:K�(%#���$nr��f?�'M����:�ǆ�a�s���~�+�r��ZO&�����M����D4��������f�~mD�%lisyx>�k8I�ў�X1��F��9#)�/(�f#"�ՒI��A��-5��X��5���ؔ��:I��Γ�=*b8!۳��L����bSߔX�/��0󖕇|�~뇆����8(3W~*�qC�S������3����[h��o�nh�=)��?D_}�K�S��Bۡ2���+V�A�5���[��W.ن����UOc �3���W �4��j������ت�$��_mW���'($g�hY��y�9��o"t����R,�u5m���l��wI��ύ�(��I�l)t�����I�H��:�ee�����q��rP$y5���>��8C!�%�,�7ְ�8P��Ke�cO���/^F�G�Uy���"�,�f�T���}������]��Im!I�������G�%UC�Ԙ �� �y1~��o�k��{2kub&�����Z�i��ZV��q.}���yC��	tP�L��� ذ�.ʼ���~�a����ӨR.�:&�~U�8W��+#e��������c`�D�2�Q�X���^we���G��:���t>h6^"�����3im� �ӷ/��D~����R;Rj�1a�wHFv��M��CC�(P��q��d��j&�Y*JP-A��A2U�����Te"�{��l�[ �:R�q�LS��-rR����s(䲴��QP#_��
^�z/�S
4��ç^�fT�&C�
b�/�@��K锋lR�yS�  �Ђ
���󔚳-}���h�\�t�cD�+�ӓ0�}O�@��8ڼq�.�o(�d�am����>�)ʙ��³	�#P�}�Ȧ]�Y�:����ԙ�P S@�i��zdk����#���qX%�+�@R����X��)}D�TֽPp��ՙ}cC0$�� �a�^�veG*�!kCu���Q�>M���-1� bº�<٬
�#��Uw�$�\E 4\�m�.p����!�P�sF2S�l��<�"��Yǔ؋�Ĉ���r֘;����$5Da�tB%j��d��=�|���I-H��*�-�n�z[D�� �Y���C�ֆE&�Z�����5�Ni��@�!pB�ZC74�z'	ϛ�*��V�T\��>�S
3�UA���
��)���Y� �am:���E6�Do�q�8l ,�i�]��a��, �ZI-	K�X��Ѵ]�y��{�U?�5�c�*/�a��Î��c	9�ir�4���(#�<�J�R���YY&B�9+�U�k�G��7�j(�r�(џ�������6�"T��+��"E��G�H����%�2HE$�7�xk���6`"o�0�[#ͺ9���2y)��0t��ʴ�Z�x����](�	������e)�e�Hl�Ʈ '��,VA
��Ϙɦ��pr �N��&�j| IP|� �C����AҸ�HR�IԵ�@��㴊^�VH��H� 3pS�/�X��r��{rr$����h�R~/a��H����\L[~5T:�'�A�JAL�ؒ�&X]Et�W���`��A;ɿ1�x� �Κi`�jŊ���{�[�U��
;�*Wu��PMGRC+ �(�p�>�
"���lT�\L�- ���%�D��n�s���\'���s��ϩSU�T5��}��+v�s�^{�9�s��? 6P���{������j4e
�� Gd��zm��tݼn�t���[@�.i)q6�0R��ܥ���	�Mم#m"�@�:+^C�xl����2!�����ma̜����J�,`,GS"��5� �\l����u��! W�\B�0�e�}"�p$���1HR�E�a�vN������H��S�o�R�A�K���d��bcЛ!��������إ�d����5,e=٫m��z\�ְ^_%��5�l-\���We�#|����O��2añz�\�
�S��p���VD��J�b;���v�u1�F5�,���J>�wi�BS�f�X��!���u�^(�U��He!�q�\�\����b�¡�߹J�m�AD����H�n4����v�Fq]��~o���6F��P�����������gMT~��螰{=�v>H{i�����{䋍��)<��/�6�d.�OCTkl�0�����g��U��}��U�Zް׌l`e����'�"��ᨅ�v�x�-\�l����#+�	����Ae���ρ�!�(Ҧ�����p���H桫;�R�nӊv��d�<�����L���+���%�XT����%?��=J�=+�<�K���I�F'�k/+�v�U��9��6?��}�Zg�*��[Q`�La�XeA;`O/V���U�;*yttȩ�q�/]!��U�"���tG��/Z ��@&BW�3��|9���Q�B_�F�-��X�Ќid�������2,O�.�!w�K�A�X]bd�Kaf#�ʀR��!�B*цQ6��q��ܴ0 t��U�A�:A�� �fcQX4�����)pH6Q���Y���y�]��i��.Ϣ��f* �nL-�v�%�]��ZMVJ����T�����l�,.LmC�,�'wQI��FS��_�8c��^Vny�Y�RL�GDAe�i5�5�W����p�0ϲ�<)̂���`��et��� 4J�><�1,	�6��)Ѐ��+>0s,���B�Y�m:AQuq��w��yV�oҎ�»i��*�`�vE0��'�ob�@����+-����"��L����H:F�_�"��mjC��\�{[�	��s=j�LG�!�BZx�z��8IՅ����.���Պ�]T��Ŭ9�ՙ��υ�}&����j��)�s��	(��UXw ��yMթ���؁μ�,i��PP���16���Za��U���X��������+���M]����(�o�pK�z_8�Z(åp�8<2��ƁұN4'{�_��)��ܒ��z��͒.�B��#S-I}��al��|�ν�

�͊��/8_�H[��.��>�,qU,��k7�3�Z��k�l�؄2�`H[�B��,k��y��T5AE@_'���I��m����	5zi��Н�Y1��3#
���<��f�F�}�;��L�����8�ź
8��C�ݑ��pz�b'���Zp���3o���[���1*����<F����-\f�}/�@εF%�Mb#� uc��}X��ݷ
�.D`5!�������G�\~�:��8�q���P�h�k5�.t�[>4��Ѣ��otR�s�	P��깎� {1���s_�,1NRY�s�ե�8���u� 3��֪����.SF���zt=�%*"v��PP�{�Ư(��5qWݼs$a�,集
,�P!��K�ّlKo����4��Y�gӧ�Wg���K����T>�3~|R~�ޫ��0�Q��XN ��˂�Gi�-97ͱ[h�U���`ߏ�j�	DY]f0>�&�XPL���\�AI�� ��|�C�|�v�Y .T�{�����[��Z�w���pж������5p��l��✹��Zs�9,r��!g|�
��7v�T�q�[H<�׀%�Giuu��PL(�TG�vY1�tn�,׶ �5w6�-1��q��~���7�n�=A���]�ɰ�%�UQL��?��ی[��������D���wcY��E7e�n�Ge��TaƲ�쮪t����:C6��J5hf�N5��@�����ӻ��j#4�5LF�wzd�w��r�Li�̭���`"�{鉱��(\ř~6T?�` ���**�V?��ĥ:�X%k q:kU�;}ͼ�Z������HS����}ZGr��!Υh�u�l�$YҬ%� �l��F�DE"���
��L.��X���@�x`�af���<�>�h����`�ff?�����A6t�^U�$
,:�e���a&x9L���bh�
��/�Ԡ��c�2���:�Y�`A�9��/��$a��硆l#n�2*�r��瞑ZX Q��QW�Y>�<�`�A�nQ�UH=Gܥ#��Q3bx�:��I���*�D��պL�����D���P�N�-��6�j�g����b\.��ws��2]�x�C�p�D�����C�G��%��pp�v^�8�yO�7��
0�la�]���!��Z��0C�x�WG�P���D�I��>��a%0��Tpa6���j:�қ���<�s/C�3��x���J�|�g�>s�΁!�C��~���}"��� u�-�)f0��`��X�1V3EH^W���Şu���ݕa��IbB��w�^�EB8��P�6ѐ��;�W�D�z��$�A72�@4Ks�z�|my�����Jn���%�����!�4!���WZ8(��iny�^�D�ZD���Yw���u����JS�� !�U"cĬ+mm�.��R	�
J
gZd��-3r
e4�4
�g�<!q���,���0�%.��dlTDd4���P����������P3�)Q�������j��������/w�F��6��?��r���b�G�%��l����`K$�I��eW�����\��7������������!�|;�>�v_���|�&.���!AA̼�l�O���%z$ϥ;L�Zv��t�V	���KQg�,�(��T
�\̾�y���~#�'�Z.[��W}6m�6�sM˻ ]
;+�@��
�}��f�9�f�G�j��1&�A���
4>�:�>�tSm�^q�B7+u��^p�mw�o��>Te�eH_5u�,^���zo�B(�bb���;����mh$�)4-�܋g�}�F�T�$*.��ۡN�W��-���,��.��Y�*v�y�\��
9��ݻ8ğ���0-����i#̓d6d�YS��Q�Q��w�43T��<-�{V�x���"DY�����OGd�q�0`�42���������Q4����ް��~������ŉU�m� ��pWDJ�ߎ٪��\U� 5:&�����T�a&i�Ҙ
/��̶���z�E�����~b4��/�E�Wg�R)_�ٛ+���5�C�7�ό�شc
�c&C�����Ǚ�6�s�U�E���2�-���aT��k(GU����'��T��F�`�o|��ȿ�Ux$3\�9&J劓����>�pn�]�	ga�1D ���9��N,��	>�8��HW��*�}�,�|�`��W�m�O�Xl��3 �bע��}�f�r���+�0�@��͊,L����{r�K2�K ��c���i1";�i����-/C�N�ZB���-9�d]Qrj�2�9N�&�H��̊���=�ϵ�4W��X+�G���0%�ݨO�{�n�v��6��#�in��$��5(
�?r���쇻H���E���1T>���Ԙ,�����6�g]!��}t������|O���Υ,�!��xJ-@5�"�*ɮ�z�+���'�S0ږ�΁½$��՛.f�3���"{C��I�B�}�>�X��ϋ��`h�ܣ��E�
�/h0�р��QXÒ,��K_�2[�>h�7�Uq�D[���l4�:�Z���ܠ�!F(�B����=����7��n��;�F����zzSvZ����fw���M���0L�T���Ȫ�#K���j�3��f��v��ڝ��wYp�G

6��c	� ��7d����^WR��2�hN͡GHC�����E0,��ʼ�US��(������5F�סU��R�)�
�X���*e�(_N�b�0f4.�>���Tm�HIIe���Нi^��M��&[���ɟך��~�\��w�Ei-��i��k���Sb�,n�<���F�sT���w��-�$�f1��s��4 �tM�Rr��b$uW����*��|��iw-���.�Ϋ�
��&��:53'�`�p2u�%#�!������ה��P���ke`�Kj�2��n����a�C��,�%�J
p�!u�W��P�$tY[U �Hw>^�cÓ������0�B�M�o�>	.�1��ݾO��!`� �1L�P�0\ڨ��r��ah�AUl"�ϒj�v�u1ִ��`=G/Z��f�����0�0��K�Q#�Q�ѓ�C��@��}:�=b��	�Y��\f+�Wt:��0�PC4좑�P4�p�Tu����,��@p͚�ϑ���a��r�n�|j�Vj^�>�X]0��T�;	]��ik����;�:�p9�xB�qu��C�'�Da�պ�0FCw�裨�������	��x%6B��ev Z�뿎Żn�x	��>tn��y��X諺U�0��ynGq����ð�I1��;o�[���Z��j�Lե�s,�9}|�C�ð�F��*�{�s�Q�j���7X������׿���[s<[<�w�󝘒3T�?�Y6�Q��� W���݊~�t��#?����)���(\8��' �b�Z���s�v�DMͤ>��3�)�q�h�5�F]��p�5�B[dՄ�zwӒ�#c�ӊqt_KTv�O��v��ۀ� 6��\O����-c<�5aF�GVm
�[�c4b�E_��W��K�ߊ>P�G��=���W�0�5��nY���Pc�I�d�k�{�]s�w5��[���'?����"��������ǩ��0+��6Q�fk���5�a�qQ��%�&8��c!�o��@	N�1I'!/W��(lyc�Q�<K���^'=68H�qA�B~���0���ep�
d�Պ%ȝ!�X>��i	�Iu	��2����G����MEgD�g�A%�L���#�b('�,?�C�x\oԔ[�%o�LfM/��g�NL$�W� o����F�F-W��A����z�P�����:�CW8��'�l��ԁ��p[��ŧ��1��,7�f>W���J��J0a��i�c0_��p�9\3h`1w2��/��X��Ɛ��!�e������G�����͉�E���\�z<��;��� Y�2L����<`3��+��+]ݴ��n�s1~Vj&���BSs�D:���� ��!��"��D{Ք���+y�ۑ�H��X�4PF��A^X'��OF�$�(���9��rNj�ɲF��^���a�,L��>sJ�\%>�6���H�Pj+~�J��-\J8��s�*�d*����!{lt���$T��d,�K�����v&�n��R�Z."�Mt?X����\^&���5bEV��H��G�T/#�ˣ�O��c<��h�m�-��lsЩ,�
|
��N}��qҞ�\V��F-�v������F�%,C)�j+���tz_�s����E��=��R�j�0S�si��l�[4��eyc?���Zv�%y����l�0i�\�Y%����p�ى��^��uW&���3����m4�Se4d��j��r��\�ء����׮���������XHá��W��9��r�3b�u�7~@ꈀ��U�s�p����i��3�z-���\�F%����Hܢ�(�W�ԹID���$0ʊ�0�Ct�*6?c6�V?jq�����䮖�ԁ��y�P{�QrG儮f5O�jy�8?����劣�cC|ٟ�/��V��u��:�YK�4���p�d������B��b�����zf���>��3�׺������h�lҠ^��f�S���*Vh��C]dj���!,,�Ccj��h�kDXL�$�z��=�Z�J[	w�K��P���]��13�p�uX8�X,���+wlP��`�Z���X�xbT�:b���a�bLD �a��'�@ֶ�z��6Xոb|wĀ'�wsfN�K�b����Q�k?�#�[��[��.�$��F�k���Z��`�#�� �O��fU�b�V����O��d��M8���H��X٢���f�J�#N��B�ZeZ���μ�"T�ieVL���Q�0��=�����D��AY%cS��A��P�S�qR��5�ﰿ�ܪ�iH�=�B��3��W��/*�͋�ُ{���oV��[�0�q'6nݩU�D�ٲu;��E�sF�Q��Ë��Cp��3l�n����a�����X�N��R��q�]D�]¶3��h�u5<��޽���_�+x���e�y�h9^f[b��p�w���}����s�05C(��QmlG_��bs�Y��Z35�����>Pv"c�����������`����'5�5k���{�`��p�����?���6�U�%.�d��G�.QwX��*��X,����{�w����;о�غ�Q�u�` ڦ֘B��]|�Y$b�(~W	}ߌS�$�50��*K�h��٬e��Cr�����2�ۮ�]����ڌj��ޔ܁ͧ��FA��p�9���5�Hs��o��G����5��3�}݀Ab-�A�2����$���G�	Z+���$#-3��:VP�1��e����p��ؼ�j�ɹ��[?�]7|��kO�G��AqMOd�dh57b4*�I2J���>����<Įͳ�=�sӗ����T,C;�Y��J��pB��R�2Nr��w��'9*��u;�VU��,�b����[����_��?v1���/��s����7݂g=���W��٭h���Q�"m3�?{��>�q�>�t��s������K.C�9����7��g0���	�ic�Қ�5E��2>��A�&j��_��C{P���/an�"��~��ֿ(d�7?��8��]hGm��]���|�tӍx��~oz�_cq� j�Z�6��uo§>�y�&��A��K�?7\w5��18���\`���5��?�J}Sr|՚-9b3@1Av�`�� �W1"7l���� ��!->|׷p�Eg���y��/�Қִ:�t��E�X.��|����g?oy�[�`�E(^����شq3Z�SZ�ڜe��H=��/�?f�؉�����'cnF��Զ# ����*|��r]'2V�DO�k���o�͠ڌ�_X@�x'���g]�{��y0���w���e�k
��n���]���/�Kq������=�T��]BF�(ǵ�݋G���q�/�<���{ދl����3P��&�����2�t�B�qJc��`�D-�`���H�:6NGX�� �q��.�K���g>K������s�t�mk�c�y��/~��睳K���DTd�%w�w�Kv����ڨ0'��?�����w�̳��\�T�2^8s�8Y{�sU��`����LqcZ���b� ُ��{p��b3�G苇��g�� ���û���Ӵ%!��}"�u�%���M
�Y"m'�V�bW�$B� ��oԞbc�� �s����P�R"m{��;w�x�ەl�k����S���%�r�
�9R]"!�r4���B6w�zأ���R�h�����g?_��y����(GG[<����#��h��Zo�,��7ߌ��/ğ��r�v`������.�o�q0���t�����(���O�g9����z����V{	ƂR8LgZ�J��$b~�0zK��P�g��x��]�L�,݃�-m���5���bt�\������'�u�����u�1.����܅�/����w-�E��"]v)�Ze��{�ޡ6G/_@%l�ݚFczڪ�
�q0��p�j���ˑ��T�kR[(敫�����()z�ƬW�<q��m$�k�����eg�Ш��s�]���06��!�i�u��WkX��Y.���L��&��A4�����P������J�(B�6i[$V�	1E8�t�be��)�q��`�E���#�*c�cܒ�5�$�CZhWW�;�f��ލ����E�,uPW$�PqA���/�u�zl<m¦�(DX���%��7��s7����/x�s18�u"7�e�aϡ�\o�μ�B�$�+y�0D��-��}# >ec��?J\9��g�UD�'Y�Ѱ��[eV�(����]���n?�n�zK["?����^�R4ڄ���h��7�WA�A������mÇ�}�d]<���m��#��;�ȽL#I����\õ�f��1�qq�b�e�Ȫ'đq�S��e#
-'�&J�a˔aHvj��g:[����}�k_����0]5\�/|�x��_����y�FYO���r�x�uZַ{�yj�Fu�N�眿��G�i���_Q��T_��7�8W�����g���v�]=��>�1�3
�Z8���:��� @俉��N~��eiQ^����p|�<��/~/{�+133��7!�E����q;�6o¥��_��c登��Ba'N;k#��m��v��>�ױ��a|�S�ö��������e(d�J+�I��G�����`gxnu#�	5�Ɏ�e���v��ߋ��r4E��[/����ϨF)~��/Ŗٍ����1,�J���n�NO�׾�5ر�\����]���ۍ١�nD�~fozǻ�ܼw��JK�Ȼ�� ��Ѫ�(`�A/�k���S��GqD�y9&k��"�j�H�4���+�'#L�7`�����;���/���z�4ds��֔�]�y�]������w�@��x�k_���J\s�wp���ik�p�G��FP��W�Vi.��_F�ލC��8�ZX�%p��0�v{�5�������\�uō���1فn�������ô���Qco�/�S����'��ϿQ]w�q'.<{7�K�8�� z����`��ͨ�ut�4��׿	O��_��7ށ3�:��y�D��0}�#EK��Ae��ulk�9x�
�D�j�����<�1t�X�I�d\�h��H�6@��j��im
�� ������c�;����o��ضm�x5�Om�:��--���o{3�x�p�m7�='�h��7s@�t�{��:bx��<	�偅:w]k@� 'S�ud�+?��p��eK`t�߭�1Ҹ��a_Q/&C7_AI���`��D��k�����x�{��v��~���Yt�0�f��3ӱ����Y�{!n�I\ӊh��s�c��qסEl:�t����	P�q��%�fS6���qJc��H:�Ө����,����f0�]�<Ksg��o|O;7�3�M�v�=�ᰂf��5���-"B$.�]`j�N��&�/��K�}K=��y�r�M�v���cv�,���xg����5�c��5����\]j����w{#eW&U����&"1,j lv�y�
9fq���;��$^���?y�><�<l&���{R&�O~�����3p��O��܅�hl�s-q���s=�l٩�}ڋ�	z\���Z��4F9ֲ˖�/�-���,�k�Ĩl6�O�Z^�����*GKv���3 ���WP,����@ܞ��{2�a"����1�s0
U+hLoD� ��c|Э�9�S��uO�3������7p������3���r�lFD�򤯋��"dX��޲i��,�gsl>�ǔc���3v*��2 ��X�{ϋ�*
�6�y�<߄F}�V�Ȉ��+\�^�XԒ�+%��/��������ʗ}�(?o�]����0��ϗ=k�3����_�&����6�1d�;2�sH���/���*Xw�~o���=�����(ĳ47���DUm�D���"�۷Ga��6�R6��&H�@N�K���+b����#l��F0�˄�V�T��KCT�R萄�2�U��A�I�	p�zc��5A-٧�Ȗ�$�F�7��n_d�:��~��ZQa�t�K4�������>��(�jJ�C�"����/�ǣ�0bT: �щ�\���ص+��D���*��ـ��H���I�����7��P�C����C�za)[�g]`�r2�d60E2IZj(��J� M�תW:���"�-��"5Ɔ����x��/�Q:�S�a�G5R8�@��=T�M�1%�y6BK��c�F�#�r�Qd]�,C>��>Eg��{�������6�/�}�����/���G��Ncl�4/�**�S����ˏ��WǄ7b�µBy�	@�b��exGUyXe$�L���=Z��]���I�Mrg,.Á�M�،�j����>��.
C�ue��|��#�+]��/�4x��j\��u4�R<;;�o�TQ�Q�D�<*Z󡛉��T�+���Mm�X		Gz�Xo�E�J��.��A4k#�q�5�֌l�)�S��ƍ;Ā��� ��FT�<�ZA���9����)[i$���/D����&5rZ�w���]FH��MA*�̣��Z���r�X��?F-��lT��zA�ץ��/�m��a,�P�_�M�D&m�hRt��V�����J�ԇ�X_�Z�X���b�|bG��x��P�Ȇr��9��W�`�T�f�`�Ar�C�؆UӟS��)*������u
`_�YZɽ��ĕO���y�]����k��M�[�Z�i��}����l�09�Z=2$�9wؖuQY}�Y�c閁���$\��f��5��O�d�G���Z�v�7�'�v
�?&�X��A*$�_�y�AODbńp������O��Kx��_߱(�p�Q���(�INdc�yi�W��rqn�E-o��D�[�LP1Ru�Yjb.�t������h�4yds��q��ɳ��e���Q��_w��tu���������e�P��5]�7��H��}��nwZ6�A;��Lz)���פ1��8��l�-7�X����UQ�Ia |�%#��%��[W�����w�H�g�`<�q�Rڬ�R:M���ڥ0U��3���v�$�i��d	?w�&�ɯ���'��h;�R���1��͡��.��9�q(����兯����(0q�x�=r(�99Y��T��UqS�*C4�yZ�-ٳE����!R[��[ɺ����}���B��[�Tɠ0H;x�/�,^�a��)Ɲb�.����Rɳ��A)�(�(C�Q�VQ8�l^����pUk.�X�?���\��1�s n���&�ŗK���h�t�f�,D�<��Ύ�J�a�:���@��N!J0�D-)�6�f3E�S�c�&�&���Xψ���������í�G��ޗRO��yZ����EV
ő¡~N8QT8\,��OP���8(I�u.�ٝ��3���P��CA�-1[�㮽�`��I�N4�Q(dÑ�%y�G��h]�@,���᠇��ѣG�e��*�M�L�b^�h�t`�C��nCv�?p�_J8]�I��t3���[������(nc0�x�K��)W�=��Z�'�����:�R��>�w\�s�>�3-�� ���t���Ck�9��[ŧ�������.<ː�s{��+�5�������� �p���D ��j,
�+RGD��5r�O$Z�P�d,��TwǎJ�kj?w<���f�zL�<�w־�Ȁ���نc�{����9d��0�o�:���hk;��:��b#M�30X����VÊ�V�Xa���jk��П@���1+36�����%����-�Xh����;�/�e��j<��y*����V������?O��<q��cœ��P�{����=yc��f|��+��>�7��qC�,�s��H�i<��+����~���ص�¯�ʯ�[�:���:���'xȣ��o���n>�#�UG�%qp�R��e
c+K����Dt���Rz1ˇ�'z�/�Y�Jǡ����!F�mPJl�J�`k�����}����'��]g?Y��D���*�E1�?�����{j�i12E�U�8q��5���,��*�w/�Z�`V���3��*�ܳZ2eZ��D
��]���V6�S̠��`wP���	m����n���,�XJ��p�Vh��(����Đ.;���O:9�bY�O��E�#N�"#5�*t�����^���)��F��"�F�C�5�YNG.�T� �P������J�(,�c�M�h�,�6�l~c�3ч�">��(I��,O2��������'��ۂ�X��o������0l�m����>�)�+[��8<�(Z���D�b?Zn~Z
�k�5��Ȯ+���G�o&��z"͙��h�b����C�s�u�Fb\�
����a�3��^�
���U�ᘞ��+˘��h���G"�5��f;�h��"��s6��\r�$@�h
��	ϣ����A#Y�^QE^o����Bc+�7
����|lj?7P������rI��J��1*;`dń���+\6־8\�y�[G��X��,�l�Ao��O!���`>�����6o�푙�Iv҈gG��Q�1��i�dRb(��AilҖK��D�9��P�b����gU��A��F2Pn����#6��6G�B�8� Oא�;��zD@�%=s����I�D,�sLM70/�e�X�$�"+Q����Y=�0�a-?�+�0��ī��q^Tk
�dN`krĈ�=����r������13<'C�f$��10��^K�w^ V
���=nΘ)F���.f[[1�9�ƝmY��y�|řh��ܠ�	���{8e��^X��dt՚�x�J��h�.Fk*��j
ݩ"@���x�6�T#��Ē�n���.
c"U��r�.A@�������@c2�#@#�/i<�F�yU��pc��-��Cr�1
k������\�%�v���&�=��#�h]�jx^s1�I/UK"������N��W��c.��e@�9 5X'��2P//��ɀXbЮ֓=I->��AqQE�'��իG�⣂̧�2h����&����r��즙Y1X���(j	�"(��l�dCl�{ZG"�K�	H~+�H�ʦB��
Y�D��������r<��eh��6:8(�l��G���|OE4G*Z�뢥�X�B�#l ��h�	R��H�~i�dnR��ж��V�3�%�s
�h5��SLe��ĖA�u���S������A��?1w�e;����QrBC�U��P�ͽ>�M��t^��	XD��\jm�0�C���O�ǣq�mP)�l���"e�������/�,l�[@�w��[��/NS�4 	�>
۸u���Ƭ�:i�Ա����%��IҤU[�z8g�n짶Hz�Rk8,�̉�PC-�Q$�<�����F#Nb?��U�X�{���b�ʭ���"�Qè��+a!L3�>�шvz���4Y�$0�&�2�Yi�JA8�`L�Q^��`Иn4���c��˼b�Ǣ�xlя��v:4�������-[eJ��p��()�?�aV�G9��8v;��	�L�ٕIĞ^�����t|ظ6n�����&�3#~��{x �;{������b;��g<N̪ȃm9���t&R��&M��/ޥj�,��f�^�|g��.A��NG��^�W��"��QPs|�EC�Ӛ~��q0Wk�QUW�8�G��}Ypf+C��(�]�F�-gwU<�@Y���⎒��L�	<���(2�Qs��=�%hb��#t�J�͗�raA4r�UU�WmY*���2Cz$�`��N�}��jr� �p.��Z�X�����8�b�{�����"-���$�h��!��vY���g�� \��?��!�N�[��J��� �L=�Bŀ:p��Y��?�!N:��qAA���E^����YK;����h�m6�_{Z1�^��x �ZZ��6W�2n�bw$�(�X��RO��b�k�"U�Ĵ�@���2��j�mlajX�,(��|��.\��de���%�V�P�3���9-ǤQ���%�F]V�#s��+��$��0S�D��Ȇ����,Z�`h�%-i�V�e��nte��D��-��]&�LŒ�ԵK�=��@]�x�A\���fԛ��W��gd�]���_��p�E�;e��C䨠��` �;�VE\�,��~����@��ކ�:��@�SC������	Y���p��h�� %�!`�
�)E�i�x��³(�,F�h4@�M��G��b�*�R�T���a�̆y��)%	�k�.����}+SQT��)�I�+��"r�����aE(� �b�����Y���xW5�™,�-�}�E�GM������yn��p,�b`���2uG���W��r�����8~�B#��4���ҵ�g+�" ���S�x��A�!�Hu٣IA�h�*6EC��"Ҙ�H[	y�e��scW�cQ�����+�ȃb�?��NTXp��b�G7U�4�IHEJ㙂�x�ުB�����!zWd��"^����(�m퓖ss�V��v�5h��p�H�s<�X�P�8�VܒO.�R扆��}��v�s�X�	wR���,�#^���S-��E�D�]�㸳G�Q�jq99��yD/D�!�4*.���q	߉�J���>H�5��w�r��5��hFa�I,��,6����Q8�\���q�VBd��zRdU�x�$o+p��Oȭ6�xc��:L�h�Ck"�$�S���Ƹ�H;1�SӚ�]�,�f��)dؽW3�|e܁@e�\�(5Tb1[U��bYeq��xz�Z�X�`��!�������$��8�1x$0��դ�Bn�(pVK�\�x��ʻ.�'A��6�=��1���A���Z��x���Z u�:��w�`��f0i�p��5 �K0\�^�����9P}�P��-�;$�6��*v��OML$Z=�~W�c��g�f/aK!G![�@'���{-�	�P�6U��rn��e�B_�q��	j���y���P�3����(B���#1�#CS�C��e�X#�h�t���o\��>J9Z1Ĝ|@*�6�ۊ���-֥�����Eq}�u᫟�\;o#�~g���/��̣-F%#�*8bwt��҇?n�X]fkD�Ϝע�:X�9=����]�>T�9#�N��'�e6�����E�u)�U&��8Tۤ��^-p�-�a��Of��A���"�zMÓ���u��Q�4�џ��M[d�&��C��w��ϽL<��z�i�6��Gj^���1ƪ������%�F�g_��~!ww�Es�K�z'����-���i�]Pm�П����p�Tf�k0;��v��X���,1��-��>KZ���U�Yո`ʅ�X��銊�dK^���5[H[&&��>���_Ʌ���(�R:��}��m�g�]��x�����/GO�d��d�����~
ؾ��6�'��K_{�֩,f^�8���dԣ�j���[O�U/�/^�2�6�@D29�?x&�?�g?�J۩�2��^�y�Lm�Q����_�_��'��h�7 �4q˾%��Wc����jaO�
T�G��5l\�����$��8�A!gK3��M3�X��7����G\����Qk��n�����n�\�+)Vy��5�ח<�I�͙a϶
j��~��E3U#��̆vY�KC�h����2N
�KK���}䪲#1�2����U�`{b=w��k+�B��[� ���Ɠ�������2�F��%i���u�#IG�G���B{%7�S�SF���B%yr�ꮲl@ٖs4*U+$�5e�f����T}��j��e�㗭Ze\a�Q�߿ҋ��%�EVVÛ��f`!���ES��H��9Y�,;���^����=���.������o�#���^��X��_)����7Y��2u�NhT�L�z�/D�����Ci�<3�GPZ�����ל��u���MvT�n�����ǆ�ѝ�Ul�l�dM;�f:�sW�r���5 g���Z6.�U�f�#K��]��xմz�aC����Ov ��x�2f��X�i�/�հ鍜�}a�e�{�uZU^�Ҽ!ih�8��J�G����c��	�����۞�o��o�uzX�R���Fk��+n(0�pƑih{�=HU�+��`<��f�'�2��D��7�B��T�pe�h��,�dWOq�C[��zR�86��j3���� ϗ.zY����.>B4�qBϑGG��*6F��-X�6��\���3B�[Ȉ��s��pe+���ɱ_}G�T|qn)%��I�����-������Ɖ
�FQ�wN����윂�D���V�[�����١s�=_�ڞۄ�s�;�q'(:#V���?V�1֮[-Wb����2ʨZ���{��S�6%��O���y��-7��+��WV��<�Iן�5�IL���;78�����z��qn�iP��լ��<w6�� 'c-�k�v_OC3��3K#>aS���
˝T5���G��u^��aBV _�� ���|p�dJ�C��]c�T0�^�ޙ}s2�K�Ń��3�%�h[�}U�c#!M��B��%���᛺���6��u+�(�	'~V�U��:�*7���=6��;�jh�G��;\�N9�8�}���7��0���bh�Q���|��sN�K��h�u�����l%YTKX�HT���(mP�:��+��݊@�D,a�Yq��F�y�(5�9������w�E�(Z��X��aeO��S�XAUo��uP�;�2��Lk跢���-v�l��e��&4���U%�?Y����Di���r�Qq�,+��,D��!���(�4�oB�r��_�_N�Z~?�/�)U7�I8� ͦ������̿-�<�k�"�]�ܮrH�YK�c�M�����(�)���e�Ga�Y�G�]��I�`��W� ��}�}��4�c��љ�<�w%5�Cd��4�����u���5�m�w��ǳ�����}v�z;�[ Ѭ���q�A������w�,L7�ǐk-�Ά��X��_#��l�(�� ��2���Ώ������P+�+)F}DVMA�Z?����ֻ��*4��i�NT�-�����0���,/���|��~��ZB�G�ח��$'uKqƃL�I�-�rN��1��(��(1�n�[y�z*YD,��r��s~W��Qva�"��h�M�ǲ�w{,�>���Q&����O^��m`��ziM༇�S�*'WY��_23Fc�Mkڊo��U`F��ベ���a2V1Ũ�E;�wؔ��Ga��^�v�Fd�&IZÜO�<`�Yl�A�>&[���� �7����Jo�w��+>�[�N �w�&�<L��������`�s-��U��"i~��!����A.G��,!]Y��΋�}��w11Q�V,�.�(\s".�MD�-=���m��d��jv�{(�й��]t��}'&j��-1��Pv���sx��������!O�
:d#U���b^��ui2�]������%,����2L{U��b���N�aZI�f��o:�_N�������c��ba)JQ�aMI���LU��L6��}�6pE�>����T�0ꃳ*e�����KP��;�X�T�βD�<*a�4�=�������>&����W.�^�%[��ܡ�X�#�*b�,��M���Qf��>��Z�jb���F�{U��Rg��+��=:r�d̪��i�v���}�C���
��+Ǒq� [���̝�'
����U���51���`��2.)�[%���Z�2Y�`1+��P��x k7iCd���o��zݎvw3�Ċv&�<܏G��I�;-�W<�������pYH���1Zǆ+6�0��j�JcF����:D'�jMk+r�īh�^��(o��>ܰ%��z�ݥv������Z�����Im�ͱ�
.mj^����la��\���̚��H���Jh�~���
ƭ�c���G)�f3�1��%pY ��u%�WLElMd2���Z�]����N.�/�5�c�����B�b�l��zl�[��!q�f��'�Y����c��E5d�����HG�?ʞa����i��q?j�]E[x^���X_�f�z�5��|�++����ވ�Y���':�6F�6�[E��EI�(tP[��U�D�S�:�y��n1ºz��e�~��p��K+�L���fD?�J���,�8�N�;;�Z��5|
VY��&�J<�td�
dD���ŝ8��]폰�{���9>+�u��AY�V�W�� Ř���}z~����.0'%�sS5Z��Gꪎ�q��C-2He���E+Vo0ޥ�$�U1�3Pau��XSd+&���4�R��ͬ�5tF�.�b�Vv�6	��T�KSm�]��z\�'��h���h
�E���r�[\��v�-6�&������Mc>֠�Q��EaU�
o���g؊}&�}�7��M(��GG�E���{ޕ�-��mP����y��cj'EiN������a��I3$���@1��tǛ��D��(��'2�$����d�5��U��E�^֘fV��F(N�h0�`Ҩ?R�B��,�Б�Ԙ9ʴ���i��H�LB�S�90ΨA)l6g>�vߎUl�����(�x@D����x�q��H��^}�@��|h;�g��(�[-�T�`XYs��D�xP��U�6�ar���!�O<��� w�"�r4vY���uВ3�a��ݪ��X�����;�&�|�f�1�F�q�s�?�fg��.Y,O��X�^^�X-W��o!�~��J�ɝj�������"�(��v��������]���6��*e���H��]�j��)G
���h���:�*��l��#�0NZ�)n����qF}�"��^����C�*�o5��ׄ@xOfbh@,�O�4ǘm-p%y6Af��k����4L~c��d��Ǉ�K�s�����e]�0��m�L�c�*��c��ǸgF�r&��~��F%6W���^g��k���C��/G��/j�k�5���f�M��ڮ6�Ѱ�Q��B����jL�+rx��
i�Mi���Q�.�gv��|������k0����������Ñ�� s���Y�8@-D��i�X��*J<���:BWk�,k��S��f��G�w0]I13a�]�����Y��k����i[q޹�cv�F\�5���7@�kϾλ���۱Y�%�-Z�1-�G���Pm������hh�r��r��������bBN��x��L����Iy%��Yۨ�	�j��qе�Du�S0�D1ĭ�� RN�I2��3���(��.w�Ot�H%��Ii	�6M��W�;������x�_~����ٴ˱z�^��$���V|������֕"YS���	;/}8n;��-;��Qo�����8��4A�q�iC�D�f%,r�I|j��ʚ�0\�D�7J��v��s�@�F�4��¥;���M8`Ho4*�����KbC]�1�[-5�r1�'
UƑH[�p!�X�V��\s����ѻ��q՛��z�c�
䣞���Y?�0=;��z�x����o����}���O�7~�٧�;8�8m*�-�0�b�����oEy�c�T��Dl����}Ѯ#ͯ����.()���_~��#���O�R����@�*b-%?��Ǎoz�|K`7��JW���Ko�����0�˞�r,UN�(n:��,76�a�y �A(F�ᥡxm�%$�Z����8��}�U��]��k?��wnr���թ��:��=d`�������?�?�����Y��F�L,�50Ԟ��:��&a!������]/8\��ڒb��a|卯uu �6;�|n�1�����bg��KQ�r��-2�H�bB1��kk��,��+������`�\����L�A#Ws�+���D����ȣ~�"saU'��v��tw��O��M�۵ �#���,�1�%�R�0�Z�T0מF֛�L��x��G���6b\=� �c_�_f����8d�����W��w��k��U���/�����Tis�ץ+�TE���@0��s�ծNe왠$���&�Ɓ�:W�}�ӱ{Ǵ�0^D,,.��`��  �:�����u�=ޅ����	��,.��,?|N4����:K'�@!������p��	`dq1���dQt��+�VbɤV�"di��S�aK�ŗ?��x؏?��P!&Vl�),�D�q���B �@ql%��ۿ�CK	���7��]��,|/]W
�}0ֆjE)��������T�Dh5�sS���X�$Y��j�1e�]mn���-.��"���K���˰�T�⚆À� �z�D�S�������+�6���d��,ʩB �F���gl�o������ܪE���Q��~�z-���(&>���!	[M�6y����|�3��~�|�s��O�|/GufZ\�B��x��d"��`y����3���R(�>;�"��W,]$.8��LOOc~~KKK�29<6�Ɏ����D+�Sf;�V��/N s���U��"@�{�^9ƕ��*!�}���1ը���V���w��� 65]<�I5lV�bJ@���G�����Ǩ�V:Ǐ~�ݯ�E>�=�hO��ngQ+��j� u��V����	-�c�!����E*\Wq&4�Yg��Zd0�(���f�]���녣�U����r�\�;vh�Dwq���H�$n,�6���w�]�y�'#ɓc^��lLo����Gr�d�{�5x�c?������Kt��0(�������2~����J��Z͚�W�B1b����ݟ�'<����A��ʱب��*�m�~���qz�y
��%��Y�R����"�B,Sn�ZՐ�Xҹ�D]aR���͊��:�_cȍ�s��W��5>�G�+b�h�'�Q�gq������v��!� ��?"�LLg�~�C��O�5Hn�F4G�i#A>��X��s�A�f�������H�!���~�9x�[���={6�G��2��r�I,��]�ڡ�J�ȴ�g?�Y\��������fu�J!��ح2<��T;��q8��v� �4;3��
9 �L���©��&�����׆;7��׾r�^0���Ƨ��SM|e��(B��G~����\��wź�UMQ9�,��	��6Ÿ��E%GV��U(	��2ţ(�;wlBk�6��zl��n�� �S�����ᅿv\�(Z�%Gk�`��H��SSSG���V��^A��v�: �D�)=��� ���X6��Wr��䓟���k~w��\Th�E����Ck'�# }'ល��O�9S�����¡��е9NqL��ۉ�:���P9�+2*�+����_w��fkZ���x��Ql��b��9���}Pkl��%ફ�£x>�h�ǜMX~F���dn�U:-��^�?��G�B��)_S�щ��s����6X�B +z���y�,;�e	����O�����Xs�ꈰ4KW��qѹ���������%Í\� 1�Xͭu�.X�W��TN���@�	�C�4��G��hvW.�ԯ'FZET�pi �0v��c�_Lj�ȴ����~R��s�?|�׷	�]Y�����]�� ���I?j�8��5�4�fx!e%:��k�������>|<��'�����Õ�������*w��U����"Sm��Ts"��ߍϊP��L4|	��y0��6$*�&]Y�ǔ��=�d8�,C�h8���0N�/��ึ������K��+~�yY��cbpM�h-���ʮ�m��4���F��6+��:�����E[�k���J����1�!(W}]N�Ĵ�ߗ='r��a��@<��n�y6�]8&te�_�n}�(ߺg��-�5�����(��&�U-VV�z�&F{����J��v0��J�ܠ�*�ipj��q�rj�D�+
l��D����PR�zlGDLۂ~�ų�AO�\���Z���+_�v����U�A�3ϣ�+�׌�`��>�[vs%�!�[u�z��~������7��O�w�d��/���<���1�Q����W��f�b��.yG���u7`���jk���MOa�)Ζ&B�+yI�ڥ��k�7y�H"~O���q�Rڷ>C�B�;f��M����;��ٳA�c�Z�i�8Q��]GW�b���v]s�r�s�N÷��C�lQa�hvO�=i��U����%��佒��~����C�B����u���B"5oU/a�ؤ:@�Gx|�T큲L8X������_�7�.����遟�.�r��VL���V���Gj�uUz�
����V^�q�E[��I��k&�F	enS3�J�=����Z�kaLIf��W�����˗���<�"-qb������i�b260�7��e�T�r������k�ť�x(~'ݭ���G���K� ��?V��e�	Q���G#wK�1M4D��9����'��߷�B��/����ԅ�vaf�z��Ny�6��5�e��� �#rC�;���P�� 8v�C&<6nj^�a����q�RBS�#�P��Ʊv���Yl����/��.��C�-�}��a	rd�� %�*�rKN�
�:T���	��S���uo}����@�ܢF0��T�r��T�
7���Ϗ�j]t�3�D3�L��4�n5,?prV���=�N�3�\�	L��iL�X���`���5�̯}�B���i�a��(߻�?~���_���k��!q��(M��f�{Y>ծ��ط <�g��e1ІU_�k|%�Kp)J`�������4��zJ�{����	���7���"�G̘D5�S���D�&=Z�a�QK�ԕ�e��!��߲��������[���������]�e�Y�%-f��n�[��;$첋��Bޗd�v��T&���/�G�����d�ғN��=뻡l�R�"��|��/�%�_��(ƅ���:��`Y��XV��h���k5,f�i�$.�]q�Ȕ~���.6o9�����َ>�����=��.6������o�lR��_��P��U*H}dB�v��`�ⓞ�Bl}�Oc�3ppd�ܲ�D���(���D�f6nV���?Q�梫��̳X�!3�r<uʌ�
�̕GM,�����S99�yX�s ���.���������蒋A����L �/ڍ��QhB���EW��NV�yB�=�]NF�2�����T��E�lۿ����E����^�
��߾NT�����5厐P�C�^�2�z�"�*����"�k�	��?~����#��Jt��R[�PQU�м���G��J�<�����\��G/:y�*K	�(���,�3�0�w��OL��o�t�����b|�w��=J�F��4����"p@��2� d�l�$V	eg���S�5Е�Ui:ɚX�����¹|&(j��/gI��P� �Bԧ6���,pѣ�����7_������YNR�{hb�c1,k>#��g�Q��[�x՛ޅ���7�G��=�OCM�)�$�C�Pu��G��k�,��KAT-X3�P�@�GvnnN4ƒv���ڼĎi /�]�6
ׂ��\�(C�c��p?���v����+��
�R,�Z-h�hX�j-��<`����$b"PRa� �I�"Z�0S�bkD0Y�^���/�S|�u���7_���b�T!b�E��}>4�j��V�/�O^�B�����|����H��1�V����u�@���ص��%䑙"&W��sG:�l�����w{%��6�T�v�T�5V�?����S���:�#��*�\w��!;���Fy�l�CY�Ly���RO�>1���� �Zؤ���#�Fz4�!Y1��.ϡ�
Nc�1:�Q��Hda�"�ڎ��<�E������az7��m��������z��
�ۋ����%������`�9x�o���v��IQ��E"�X�A�K�lP���!�C8��*��`Q!�蛲��Fg]�����P���nʤ��\��{�Ur������Z��f�20��&� ϱ�aB;첱<)�	�յ�-TV�*'k�7.u�|F�?��~���)=;ϊ)<���ɉ�]��F0�"�T��dd�!�HH΅��`���~?�x�q6�x�ȿ�7�x6�����`�i�7ƕZQ,�o]{>��k�;��
8l��p�C�{S{5Y���w_c8�g%܂�Q�Z���"涊��xdvI���'ی�,q���B&�R�,,P�ƐH�]�j!�Ո(�#��ȵ8�e`l6��']��+��8�.�RXUKк�X�ьR���Ri�j��-�"gdC�}�mŰ����k탇(�G�4S�E�eYZ�f����[ο[K��;o����x�k� 3*������Q��坿o����z��6Av�p㐣�	�F�11���L�3�9��xt�8��!c4g��8A\ Q@Y�fiZ��n���������<��}�{o�UTwu���)�����}��>�������Y�S6�$��'7?�=[�Q��n<��@�V���[�K�#:�����X�.:��U��W��V��Z3]y�����r�)1L�}��F�y�ݻ��k���UW����/)x��d�u%�-�j2�8�/�����m|��FB�C��O���9'r+�Я��gj�;�뱃���	����b�1�������/����1�-��Y��Q���*�l<��߉���S����ִ�҅�ƙo�0���7/�Щf�hh�X�s� �tUL=�#D�n��C�
9@SعR�8eۖ�"�g+�
n����_Q��9����&6]'A�-i`�QIٜ�1�K VYr���L�1m�&Y����O�"�%Gp��,�
���|�T��b�`"<���B1�y��@|!�V��vӱ-����V򒁉 koK�MOs1e2�`GC����K��d�S-R���S�qj����s_KۏW���r��Z��o�a/6�� �<wi~'��71����<�M"��
�JϤ-=�>#�v׫"m�X���|7#Y N���,�(�\-}n���	�DcV�R�`�Lf-�r>5��٘E�O�3SYe�FE[�C~r`���,�?�h�\�˼2�fc��v�1e��z��(J�J�kk�P,Y~�,���
�;��{�4)��/�5��cU�2����b��yM�Z�G�{���C�X�Q7%�.������l��-C�kj�=�^�L-h�-�b�pS��4NҾ5���e^��⏃���1m�8�������tn�
�1�.?,(>�5�S�ȹ_�M`��g;yߴ������b����l
�1Q�߬%cA�e�kMy�Ai�vD&�cx�J��-Y�mtd�X"I�E���x9C���&Β�OC�g��
Lr�q��5�{�հ� bh~	5b�,����H����	Ѧ���b%�ܻm9_O���!d��@��Bƒ�J�f69Y��U�4�
�K$Mc�6-�+��s�֢�U��6���t}�7ѥ�S^�d�X�}�z�6`�َ�	L5yv������\�/;�b����-up��r3������	�Y���B*JS������#!MS?��%�Li:����3iS��&Qm�jV���B�3�vC��3JF�A�p�k�.���h�c�v�L�u��%�,�����T��!&@�31O�l;��a�)�.�>ĝ�:jrjU7��e�l���� 7���+��a���o�
8�*��9G�A�RR�����rt'J{���MN�5��d�#6�ݜ��\a�d�D,�oX��;&I���3g���|>Y ����b�R�W�ТN���|[A�V
d��V�Հ[�+���u�Z2�Cc��:-(�؆�^j�����P3ju7;��6�u��!�ԄWC3a7A���0y�s��	U�0�N2�EExZ�s�����v�VdbҮuqX�{E�|�oh ��CՕp�	&5Q�X��e�f~��U'��z���`
����C�,��g:� �5���{�&��Ս�5��&,bm�h��h%�*)lH߰r��]���\�G��y�ͭ.�\��:�x*�sZO��vsm�@�+j���� �3ϓ�|8�Ψ�E=Nlu��mi��,�ew�|Q����r�)�A�W���%	��+'���k�Y1���]��
=�]�MPP�2�'���H�$���Eiw�Ԃ>hT3	�e7Α]X~f"�f��R
;���H�K^`��.��EK�ƒo��d�99*f��
�Ŭd����&���S-~f��XJ��)�f���Z(����y�٘yNgi��&��{�\ܥ�%	'��_|����ر��^)h;�o�P ITS"�Q��Nd�+MA�X$���b�,xWI��]C&� ����6�����{p��g��֨��/U�5�s���3�����q�a �-v�)}c��5_S;#*�}^4aQi��鉐6Zu�Dk����h���B��<�>��M��T���+rltŪ1����QI@�YO�H�S�/yH�eX�wԖgU$�<��;������d־�\��W�c�J�N�&bKw#���^8�5XV��yY��� �cS��P.�B4B�1d�\�2�RK��I��GP7Mz;�#���G���xg��4���Y*:&�T�B��&})���,'�MY�xj�b����x�ٽ���T��^�Xhf��d磂h���aW��]��y�0��F�#��"�%����a��5Q�IꚲG򋤖��H�%	wD�1������W��b�T[y_"��Si��B���٢���!C��G�g���*ʎ���F�HSi�S���MZ>(����ڬ&_�\6�c֓�4�'GFsF�rX^'�$bW[����N�7�7}�أ�:T.�Y�5	.)��/��7ɸ/bkfy��!,V"ylcnF����kI��`;09n�r�����,(�ʂ��y4��-WV��/��r�䰜"ir`����,�.��9&�����Z_�h2L�6z�&�`��;��P����U1�`��VPk����#aH!''psr�+^ ���9���rbB7gw��U��;6�QW��ب��j��ۗy!CEu�T�33"�r֋�*��k��&����햇ju\ k���1�����/�!y��'�]��T�sZ]y���VQ��\��}�w=fL�[az9Vrh�Mc�%��ИhCu����(:��%���"��u?0AE�x&�M��=���:�
9N�{p��c8�����0|�i���-���<�\l}�)1	c�h�݁sљز�Q�|�|P	�e2j��a��2���� ���5�#��k
�a{W0E�1"��W���k�И�����ĝ�������Gy[f"�ΎB�w�F����ry�蔕(��("X�>���{��`���t��L�,)�;1ʲ�W!��Ƿ�<6!�{��?N<q��.��8�����W����/���-pE �����q�Y���'�C�<���"L�\ds8�2R?Y��XL]����"���)z=�eQ����L�8��g��W����gw��t
.�����(�[������_(��)yE=���k���k��O\��\v��j���D��t��Gb�Ƚ�2��;d�����k�;	����������F���������^�w��7��~��r�;X7���{���{p�+���W��ct����+�a�N��f�&Wk3�~�p��+RS�없Dc4�r���~u�����K��{o�[�r%���3����%B��޻Lͅ��!���YGs��5o&��o
�'��ʳOö;͙��a	#u��h�Q&�TZѶ��M�1ˡkhG�J�d��1���P|����ӂ��������o_{>���?Fm�p�ӣ�n�S!�>4����?˱*��=�c�����m?��-�&&�+�1�u~م�}Er��D[��;�߀��0���"�I�"��B��.������L�;��s��-�:�����!f��{�O�Dy���ˏ�	�굸�~w�8(J�!|����g&����v\��w���l�	ڙ¥g��~�;�\p��w��ߠ��l��s��1��k~�
����}��(.��;V1G���.$QgqGփ`��M�D��y�u�Ȅ5j5��qf�8|j��ȏ��^DZO<��%��wn����>Q��h$f��\��	/74�6[CT}�+���(&6���^3��*:/Ml+q�����σ(����+O��:'���~��9�:���ߎO|�2|��7�L5߸ �07ׄ@̱6u|��:�k�|�F\��Y�M}b�E�g���$��Π$�xσ��o��ٯ�ת�������w���;n=�Qǋ(�R4���U��tF'��\���rΠ�Bn�Q��:/�����]w����β���׏�=덣�W�O㸕�䬔�#��[�S<���8���_�"�H���-y�zm�6[*!����ΐ�jc�R0)�ֵ�v�Gan���D_�,�˱t��S��xIP�`���q�
�:���߉�U���Wn�����������D�4�z�E�4��T�ڢ��N�Pm�ͅI0I�&���#|5<�Z�Q����������.y5zH �h��a`�����ȕjJ�ҳYKIN�Ǟކ�_�U���7q�2fĢ��E^/i8N|�\���,����<�� ���y6�����j;vlǘ�m�=M4��q�ƺNǴ!�ã&�W^7gń��l����<*��J�*�OU�擺Y�p���73!]��O`V���Ę�B�%���7ނ�Gc���R�c����0Z^�����߻_���`ƟϠ]$O$�Q�+�=L�މ�+����4�W�*���FPA^ݖuuOn�!��\��a�9����w��:��ΚXh���v����ג�[y�Xe9L���E`b:��RQcIGb,�%Nn=��X���[(���"�ڻ�ֹ8�k�u�n��|5pꩯŽ��BvbGk'�]�m[6c�3L��p��ER��KLy��Zr���u�8�4tF?���X�UJ����b�ú��bӶ]芠޽���J���VKZ%����v��ǛE��
8&&�"���|^�g�h�����q�[~�ݹ˦��"u�%=6@��v~35������;��4�7=���j5yt��wc�Np�l-��gZTc���o^��7�{����X�Z0�Zq�H�\��xP_�Xr�Ĵ��m�,��a�7%�r<&f�f��L�?�p���l3�Yg�ؽ��!^�oz��}'`�ګ�G,�+.��>�"�>|9N���e�0GrX�k�i����Z�ZH��t�n	���؃�}�
��0�v�Jƕ>�NΥ�	f�9Y����u_��?��I&�g9�¹��A]>�����o�����;Q�2b�#u�G�֘�1+G�H\�T��b~7�|>��_·nK46N
��]�㲋�����n��j/��W��y�w��O\���x+yR4�tξw��\���%\�\�Șah
�֓��6BKH�J�,z�����|6?��y��V��A�����<��^��?݅��;kN�㺯��]�?
�z�L�|� �;�߅�b�TG&ЊM!�U��N
�ɍd�c|r~p�#��&�]y�&��]�ɗ��^�-�o����L 	J(M��O}�Q�Ys<vEں{�z�$������	<��^�i��V�1���em��h��h����Mw��-<���P[G�-�?���pʩ'�7 ��~��=�1���?�c�uڙ8���`/1oxRۓ�z~+J�1,�^X�8�Y)_�c�0�����J�7[������U�}���Ҡ
�6nA�H�}�I��ûerD]�{<Y�T&��z�V�{�"Z"��<}�����N�yL2-�X�t#Gf����t�FmǊC��ZA��06=�F�m���y��&�{�!�6b�����>�r�iN4LՕ'
0���P��N/��61���c��0��Ąn������ڔ7j��ʽtEM<�m/���S�L!V�	�� (O`J��]?} w���L;�ȊI89G�[���s�a�B�n��b���J=�.*�5��07�f�&�Lݣ�95I������SutR��YdS��Y���4�b�QlZy���8x�X]�ZH�E����f�V��� M�_!3�=�Ֆ�ntM9�b`�R����{O���k�e�6�aƕ��[BI*5yF�¸��W�8��mkg$Zn�$���wCK��_�Gb�n�BQ*�I6�6�r~(����n�����8>����2Bȸ���TC�j�m���fՙ,�/�P�%��[��$Yu_A$���j��9e5z��:���lƒ��<p0�O�g���fFj}v�����hn�>r�os:L�j ,�,#�VEw~���S7�8��s1XRijK�L��.��[(��+�6���8�9I��+Ô�P����@��*�дgBNfڇ�R*[�]	�ѫ+IM	�YN��k�H̸dȘD��A�f�w`��v;�?D&}/���6|�,1]1m+%��wuA�W��>��,:� �.�9r%���P��"*xn�/0ĲH�%�i����3YעB���1�"_Y/X�i-ñ���Nb�gW+�px4:ME:i��r�C�%�]�ˑR�g����4-k�|6���AH�� MFnv����L'1�_o5ܒ�0^��q�E�1̙��>����%�D X�����m,??���n�G1/��4�5��}�}���[��(�=���0��~ـ����I�Ք:h�<jXGܙ��_�N��=�S=6`cv�y>���{�s�[�����g�M���Y�L�C���Z�GuxT3��-:bAl�n4�I�T��w�ƈzi�� 2ZG�3FA�^]�����_Y#k_���Y��K��Bh�E%�d�%˲���~��k����U�@�ڲh�bT��G2�)CLb;�?��ɩŶ�,�~i<3V���|��	5�[�N��~��:�X <2��,\ʉ�x2��vD>�P�F<��M��^̳F��l�'X�7�XԀ�G��K��YMg��؆S3�dwT�t���|�������}��2{� ��^��J�wy�PALu&�v�Y��ǒ��,�a�t��J�����f�h��ҋ�9�\D3��i󖬒l@�M�`
۪UK����/�ݬ�Yi��l�T�~��lz��m:T�k5�,�\�[�[�i�X�	��y�ġD��L_��L&��TL��M��fǓ&A��ep=��\7�f��$j7�a�Sd�Q�PP�D$$E�m���C����󥏃���1�ť���c֏r"S�?���5�f[i�>;0˫c��E���O��n�8����3� K��h�2��Dq����[�J3h��.8Øb߮:�l����P��hE[�0Ɏ��T���5�A0�\�J~_Mc3����J*3�=����Ũ�v���Psj�\�T�Y'jj��tvvZ��e�Y�+�0$p��.c,�����݁ߘ���R�BFJ�M�S��I-m�vc��u��j�|l�8��i�]*U�7baP�n�,VÑ]W�(��:äh�h'�����I\[39�HLN��&GՋ\<ϵ)�L��h���	]�^�B�ߑ���g����#U$Z����=�1C��Sj�����g�7�I=F/����� s5us�����"�֎��쎒PkRY�C"�?��ۊ�]m�j&��x��<�Y�K�+:U���k�t��f�f��,C��5���c�%L�%���Tr�^ʤ�G'He����v��R{�� c#Qqj��z��w��ۨ�b�G�I7����`�E��8�'aI(�t�~�i����1��uy�jf�.���jO[f�����D�܍Z�wш�9����~Cch�]��fn�5�Pt�&�DU{����/�FzS�jo_�s�xz��tP��Ư�g�!���j��p��?�-O>e�J���e�%�ݘ�1��4�3�d���Z��\DzL2�~���$��a�Y\��s�n|�~�j�l��Ŗ���0��B�%�ϬtP�{te�eT^�bM(ܱS�����SN�\'���$J�1l+δۄ��4=]t���B��	�X�UC,&��f{�+VL`�ʕ(TC%Jcy`�e"������ڂ9���V�1��;�Be���W��>
f���n��L�g�Zt�E�C�d��I�Z�Ƥ��zH��q��VKwp�
�U{f"�l�TK��0u{�ڤ�1j��hʢT��-|25nd-�)��U��wH��1?0�5��G�O�n��<׀�N�!ɉ��P��R!w�[�$�J���!��APNv����Z�S��	v*��FC�ZM�����[��<l�!A�K#�9,<��A�M�7Z���o��p�f�W�>��
Z�϶��rrg ��)=�CH��}�J�{B��s��'iڗM�jm>�(�M��e掺I���	��YE���ؚ٬՞�<K|;}W׿�wA�"��Ts�m�=ǦO:�ݲ���B�S��jwǦ⩊�S� �-��p,ڎ`�PS���L*;�\Em}v,�r����N��_�l�Z� �g������ɤ�ϜI�`�g�zb,&�Ȗ���v���G2�ˬ�h@S��3<���1�*Y2S�Q�iE΀X��Ƭ�����hu{~�Á2<o!�J�@��]���=�6�<ƞɈlNbx*L�(GU)���Sx�hV��v_���a�}��n���ps�0K%����K�kL>�)2��*�%bIP�źP>V���׷�%��d�Y}��\���U.>���YI���j5EӸ�T�U�`9fU~��'8i��4ѡ5e��quc��D���$Y�Q��f����4�~^F=f�˘m� ��1�	���`Ǟ��9L�U�]M��,SW�)m`�bH�*�}z��2�s�d8����KQ|��U��٨��R�\*��@�VIg�"���)���xP&Z�`�I�Q�X޳���S�@��ݘ�������A��C�=�m:��i�����g]�f$ڔt�8gI�.�(a�gԣht���he(��j
z��,S����������ʨ'��MicS�d"Q���A1fيI�P��pkʱY��H�-dHk"�Qά���f�i�bF{e�:�b�ٽ����1��Z���O~.��mHfg�b��"[7c�.R4t�PvB�S���gFN,���4��FMP&�K
��{��4r�u��{�9�t�qfy}qT�gO�56|����~g>�g�����=���
��bQn�>�@�'�t�5�fo6��o�Y�)�\s�k�m�d ��G��f )`B���S���ȏ
���=�B��i��a"�@�0--w)IV�jg��0��3-4Km�je=B���d^[	Oש�B�u�NS�V��
Y]�$0�����ޖ����2�$0:r#�Ly��b�fy���p�H�e=�M��3t�Y� �D6Dq��
�m�HyRR�Fj�����ܘV�i�΁����P�ˏ��t�m	�����)���!i�l9H��OTS�-�Z����I���+5�:cΣ�.Q�����NK&�.�2��_��+�{�pjd��[��\�<fe#EE>��06���רFI��@vl��x~>�D }8�y>'���b�_������J_�fTE ���$,������Q]�mnik�x5�g�@ǩjL�����S�F�l�+j�԰�e~�����*�[Q���\D�*������{�pN�4�:ن<��X��.�U��@,'1��b�9%�˫А��jH�|�Y�c���g��� G��`��t3�4_�$�4�i�D3M�}%�=��E�@D�1fs�����	ztݢ��rSC���RfB�D d��_�
x�����j�tt�o��;��m,]o>6�GY����x,�NytT�挋5|m���pJU�Ϻ�cȻ��E�p�Eb%lD�Qv�f;%��2�8�o)��9���N�xEF6Mb:�XFY�܀����9;���Q��M8$J���&|��;�"��l�*�\���Z~�d��d�A���1�;����_�����j]�p.��e,'����Q��I�I���D)[)�4/�-:2�,��r�Y"V���7,s"�*�zu���� 8���u%{N�k�
�d��'M�O��f&����۠)Hb�VB�9�T�ihW�*h�A�(���ޥ֘�?���$�+0�6!/!���`w欦�65�ɓ�yyͼɵ�^(�/C*|Ij2�� d���u���NL��TK�r��Ӂl$�.�3���0f�%�R�JD�%���s0&���G`�,��؀%�z&3o#G�5�-�:(��+g��/+/k/�'�0ǡ(�f^�C����k�(w=8��7�'��Kר��-��p�Zu+k��t"s�U��O�AG@n>ߑ�5���"��vC��	��0A&(1�SqR�������f��O6�Y�T�+�u���ԛ@�SG�K����䞺ih�H�^W⩮�0W혓�(X�A���`�.8�RDCE6M�`�]�-^�G�rd:6�L�w�ɵ檓�I2_ej�2�s�r�5��h�S+�y*0C��ɤ���b��b��Uu�%a����[�=E�u�[�9����u c8j���cCs4���|�/��#�8$d�]4SB����=�;m�}B�{�N�i�`�+���Hh8��	4��8�<�иè�e�ш-���X7��	-'�̙�Yģ�ڋͳK��Ԉ�蘒��`Q�}���ibx�X	mG1	���E^o���3�Q�T:�}��"['��,�����Q�nhh��:�M�I@�fV�(��\��ȘoZ��(�{��q]ߓ#�����6�v����5�FNO(H����b���z"���Wa$ECО��B�]��X)��2�<�ג�9����O3�f7҉ɸS=]k"g�+M���?��S��(3a$Z����d�b����	f{�q'	�'uc�IO��H9@�U���J��.`d	�����O�V&b1@�s�`tc�\7�ϹCb�9i�T�Փ�CS�x�ߡh��Wn^�"Q��y?�Ė/jy�Q��p�-TGdG5v��D���f�i�b�;���9Vx�DF!���5NJDǸߍ��|�:��sI.g�.�0B��F��]Y�Ey�1�gŁ��j<�q��0����h��>�h̲mu�K�����{�%��A�a��e��1���T�݊�ĵj��YBN{'	،v� 	��ߗ�):�޿c��C���׼t^��r<G= ����~�|�=��m�[��"�yG�۠�.�Fԏga �!���W=��:k��� ��Ҵi�E�p.�̟x�BŐ��ۋ�ʊ������H� I㚝h�b#�^'�B��=O��@OuQҸ�=H��5�����������S�v����Ǣt
�>Wұ�fKE��g�G=���C��Tk0�<���v|�ǳ�Ug|��z�0�[q���\vT>�|Of�4~��|+V3��h1�Ӗ�Ԛ����
�o�ƻ7�MC�9\ks3N�&?��������a�El�LD����az�?�隴��/��;�FF�l6���O����?�p]o�k;w<�X�Vav��7O�����-��M���շ�cc��x�ٍ#pm���6�s�|�������_L��%�\	�\��_�η�������������߽`>Ƶ���^��7,w�,������۱�T������9�\p�,�а��r���߿�'����ј]h+���^�����6��f�v}����N��/�(�l�Y�c9��P�0�(��8��_��:Ђ�a�S]�k�A9�ꄫ
��rX��2/?����A��D�B�GqS����Ǳ��)�1Q��e�x��I	,B�l�Q����c�ޘ(V�rf7��/F6��wʬ���֬Amz�����n{E��n�y��W�57s<�q�K�D�^�Hշ��q�qL	F�T^YL;�3�U2����ɏ_��|w(_*�_��bg�b�8�4ʗ
y��d�/�(�cJ0:����8��b���0q\vC�>�sD�'�v$ʣ�>����e{�cJ0d��O��xK'�\�p�z��ue�JQ��'ը��7��q�	�<��4M�M0r�eJ���/����a��A��˭��֣z�k�����Gl$��KO�^�؟�`���8�#]47�aG{.�0KGq�ɘ7D�� ?�C�����R1����O?�`��w�r.�����V����hjO�G���ڗ��Xf�8��_�c �l� ;vY����L	�Qǔ`�_i����r^�c�1��U20����5�����܂1o-^��c�s}�Dq/}$Ird,|��_��1O0�Y��s]�h/����e�d`̋O,��V�����Q�,�bj�Ʋ�ǔ`d~Vl��5�?D�Aļ&��I��|�M������Q���.'���(��m3�	�V����jy�Ϝ#��.�qL	F�[fa��o��,H��lCCCڈ��l.[ȟ�����5���pS�Q(��Z�P4E�NҞ庶��z��Uv�zY��-��2��cC�,��]�V��Qǔ`\|�ş���V��eq��1{�r]���/���۷�#BY��7��n,���K�X���T�3r�8���6�o����q�eU���8Jc�ڵO�ǔ`d�h��c��W���3j�    IEND�B`�PK   6}�XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   ���X��N�
  m     jsons/user_defined.json�\�n�8~Ç� ��ߤ�_6�ťI�����"�VXG��v��b�^��(ۉ�d���l�4��oF���p�Q/>����x9��/�Vuc�x2�h�y�6�8�S�̗e�||�����m�qg�uӎޞ_��Z��m�ٝ8~]��m�����v�������Q�fs;���1&�d �@P�����$�`�R�����uW�-�Nn�_��}�(62��@2#��[M1�JL���귲GP�{8R��eӺ/���US�������������v6�}-�̝�=~�ޯ�����QZ6�oK�Q��\/�ڙs�ٟ��������A��	��������]2>ZtK743U�����o�_�����a���a7C�������?��x˒`���.��d˓`ɔ���!�HBeaL6ĔI�/���A�g��(�I��ܱ���$�c�,��<�Da�e����àCQ�4��0�PR8���4:N��1��Tp��A�O�¨E�D���0�GS(�8 �PV���Ċ��B$�E�5����a!`O�b��a�bO�⩰���=IK$�aTOΒ��2�:��*j���0�Pc%��0�Pb�d���2ؓ�H"j8 bO⢉�ayaO�b��auO�≨aqO���N[7�i�ump_wn�����M��l�	��`�%��Y�������
+�!�f�}׵w�[ԛ�aSo�׎�9�����k��C͖���y	yO8wo���C{ќ��w���Ļz^�3�x���-W��&����,�fY)�Xv�0�1�.��i7��]�6�Y�{����[�ޞ��NZ/3������z���Uݍ涙���Im��y0z��n6ET�vǁ0� �
��K���r���~�Uf��#�ؒ�c���[�tŖ���V�Z˔��lÅ-��ưB f(�c���\
fK��.��W�L�S7\�*5$��q���0�S�9���B�UҍTn�2\EJ��П��}c(����Q�P4��Mfnfnfnfnf��܋��#��'NG����u۴�C�����Y�ޝ���6�g��rq����zXW4�HW%�i�	T�P�&\0b�+jR�g��%��*�t��$����VDR�	���[HΔ6T��=}(w?&�T/�}6}ݳ�(����;����/�hʐ�;)d1e� _ �{H�����1���8�a�_�d�����>��t�~-(E"޸;ԍ�����};r�F�����2�!)$�$h�©csha40�0�[+�ղd��67�'�I�Hŀ�\���*YP�R���i��������/T���}<���[8�ˮ�,ۘ�9�P4�����'�����Q{|A�Puf{R؛'|Q�ʙ��g/g�\�
�N�0p�˳���ꋾ�LK�l�����O��'�8�3*ܳ���m�۝��j�t��?�X沃&�*��$�����~��8�5�5�5�5�5�5�5�5�5��/+�׭Y�����*i�RD�VJKJ��
�%**�x�W+K����L	� �ZX �-,J)),�(�9-�%���!�(U@�

ͤp����1E�b�r����{Gh�
(�AJ��U�Gl����澭�"����2����A�~��"��"/��	$/���/翸�$xD����y
w+�x!$�H1ܙK<�*�J+����x�����P[��(`t)����M�!VBs��0����1�nb��"�@i�p~���w^����rĸ��O1D���y=�#6�.,�	qT@����i�[-�OC����H#P� K4��;�<m�[<�@�?ʓ^��8��,���H��7~Ğ��-�L�7��ZT��'���4�n �l!ܱ��[ݱ�R-D���,B�4z�½��v�]�X10nB�4��H���h�@�G��������"w�4J������Q��q����Q��q�c<�m����<]����yE�ӝ��OU���Hu�i�凧�H_����S�u���Ӽ�5���#/�����)4V�zZ���94�������D#-�Fw~xő�O�;?<���+ 1)�'Q���f��s(	S���O�$���sz%�Q��99��$a��������y�@L�����2l &����"r1A'gN�.Bա������.=\�y=_�ݓe�����k��T� H� �)�+�)Zj�Ʃ=��(�8-9�JPr.0$���z�$��/z�@x��2a�����H��|�̄�����eO�0�����>����A;=�]��?�����`���N��3��kY��������\�潻�g8�����6�qΘ���~��l�ow̾s��z��p�W������>�~����G�]Ot�~Pp�i��������3���v�6�I����$х-���oa��h	!.�L)��>S�9"䈐#B�9"䈐#B�9"䈐#B�9"䈐#BjDpn�:�P@���I�4��[E���c���Q�%�cX��Bb��!��L�b�-,�4��e%*3l(wܾ\ńMS�Lu����5�(��5y; <[�O�Q�~}��гZ�:Z�#k�Eߌ��W��ѿGC;G6�zϣ��OuT�껓����^|�|��E;.lM�J���k��q�������?W���xq���M����xB�APU�,�����bǑ�v��N���>�̞�qɹA[9NS�-сDBR�a%ʬ���������������������翔�o��PK
   ���X����.  `_                  cirkitFile.jsonPK
   �{�X@��)  /             /  images/0931d3d0-b3b5-4a2f-bea7-013f7f069bf2.pngPK
   �{�Xǐ]zd� K� /             �E images/0ceeee3a-ea03-4589-bdea-2202a7c6e233.pngPK
   ���X����7  �  /             F� images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   6}�X~��k�6 4 /             �� images/663b53f5-e86a-4272-a51e-f5b809259b46.pngPK
   .��Xd��  �   /             �	 images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   �z�X�ة� � /             �5	 images/8e621aff-3cab-4d84-92e8-90ee5aaf6d75.pngPK
   ���X�&�}[  y`  /             �O
 images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   �z�X�H2�    /             k�
 images/9865acd8-fab0-4625-b565-b7238dff6b6e.pngPK
   }�X��$W� >� /             ��
 images/a4664b0c-b4f7-4551-a44a-c7f07c5873cd.pngPK
   .��X	��#u } /             o� images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   �z�Xk���  ��  /             � images/aa6b0e15-4878-4df8-8b7e-ef384cc3161e.pngPK
   }�X�F��^ ~% /             �� images/b0a0d881-65db-4735-bc7e-86e9309b8843.pngPK
   6}�X$7h�!  �!  /             b� images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   6}�X���]  [  /             � images/cbec1558-c992-4de5-91c3-4ac90e5ffec0.pngPK
   �z�X��/F��  ��  /             � images/d4cdd597-5d42-4626-88f7-26875eb62832.pngPK
   6}�XP��/�  ǽ  /             � images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   ���X��N�
  m               J� jsons/user_defined.jsonPK      R  F�   